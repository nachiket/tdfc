// Verilog inter-page non-input queue module for JPEG_dec_d1_ScOrEtMp0
// Emitted by ../../../tdfc version 1.160, Mon Aug 24 17:52:43 2009

`include "Q_wire.v"
`include "Q_wire.v"

module JPEG_dec_d1_ScOrEtMp0_q (clock, reset, outA_qin_d, outA_qin_e, outA_qin_v, outA_qin_b, outA_qout_d, outA_qout_e, outA_qout_v, outA_qout_b, outB_qin_d, outB_qin_e, outB_qin_v, outB_qin_b, outB_qout_d, outB_qout_e, outB_qout_v, outB_qout_b, outC_qin_d, outC_qin_e, outC_qin_v, outC_qin_b, outC_qout_d, outC_qout_e, outC_qout_v, outC_qout_b, outD_qin_d, outD_qin_e, outD_qin_v, outD_qin_b, outD_qout_d, outD_qout_e, outD_qout_v, outD_qout_b, outE_qin_d, outE_qin_e, outE_qin_v, outE_qin_b, outE_qout_d, outE_qout_e, outE_qout_v, outE_qout_b, outF_qin_d, outF_qin_e, outF_qin_v, outF_qin_b, outF_qout_d, outF_qout_e, outF_qout_v, outF_qout_b, outG_qin_d, outG_qin_e, outG_qin_v, outG_qin_b, outG_qout_d, outG_qout_e, outG_qout_v, outG_qout_b, outH_qin_d, outH_qin_e, outH_qin_v, outH_qin_b, outH_qout_d, outH_qout_e, outH_qout_v, outH_qout_b, ScOrEtMp1_qin_d, ScOrEtMp1_qin_e, ScOrEtMp1_qin_v, ScOrEtMp1_qin_b, ScOrEtMp1_qout_d, ScOrEtMp1_qout_e, ScOrEtMp1_qout_v, ScOrEtMp1_qout_b, ScOrEtMp2_qin_d, ScOrEtMp2_qin_e, ScOrEtMp2_qin_v, ScOrEtMp2_qin_b, ScOrEtMp2_qout_d, ScOrEtMp2_qout_e, ScOrEtMp2_qout_v, ScOrEtMp2_qout_b, ScOrEtMp3_qin_d, ScOrEtMp3_qin_e, ScOrEtMp3_qin_v, ScOrEtMp3_qin_b, ScOrEtMp3_qout_d, ScOrEtMp3_qout_e, ScOrEtMp3_qout_v, ScOrEtMp3_qout_b, ScOrEtMp4_qin_d, ScOrEtMp4_qin_e, ScOrEtMp4_qin_v, ScOrEtMp4_qin_b, ScOrEtMp4_qout_d, ScOrEtMp4_qout_e, ScOrEtMp4_qout_v, ScOrEtMp4_qout_b, ScOrEtMp5_qin_d, ScOrEtMp5_qin_e, ScOrEtMp5_qin_v, ScOrEtMp5_qin_b, ScOrEtMp5_qout_d, ScOrEtMp5_qout_e, ScOrEtMp5_qout_v, ScOrEtMp5_qout_b, ScOrEtMp6_qin_d, ScOrEtMp6_qin_e, ScOrEtMp6_qin_v, ScOrEtMp6_qin_b, ScOrEtMp6_qout_d, ScOrEtMp6_qout_e, ScOrEtMp6_qout_v, ScOrEtMp6_qout_b, ScOrEtMp7_qin_d, ScOrEtMp7_qin_e, ScOrEtMp7_qin_v, ScOrEtMp7_qin_b, ScOrEtMp7_qout_d, ScOrEtMp7_qout_e, ScOrEtMp7_qout_v, ScOrEtMp7_qout_b, ScOrEtMp8_qin_d, ScOrEtMp8_qin_e, ScOrEtMp8_qin_v, ScOrEtMp8_qin_b, ScOrEtMp8_qout_d, ScOrEtMp8_qout_e, ScOrEtMp8_qout_v, ScOrEtMp8_qout_b, ScOrEtMp9_qin_d, ScOrEtMp9_qin_e, ScOrEtMp9_qin_v, ScOrEtMp9_qin_b, ScOrEtMp9_qout_d, ScOrEtMp9_qout_e, ScOrEtMp9_qout_v, ScOrEtMp9_qout_b, ScOrEtMp10_qin_d, ScOrEtMp10_qin_e, ScOrEtMp10_qin_v, ScOrEtMp10_qin_b, ScOrEtMp10_qout_d, ScOrEtMp10_qout_e, ScOrEtMp10_qout_v, ScOrEtMp10_qout_b, ScOrEtMp11_qin_d, ScOrEtMp11_qin_e, ScOrEtMp11_qin_v, ScOrEtMp11_qin_b, ScOrEtMp11_qout_d, ScOrEtMp11_qout_e, ScOrEtMp11_qout_v, ScOrEtMp11_qout_b, ScOrEtMp12_qin_d, ScOrEtMp12_qin_e, ScOrEtMp12_qin_v, ScOrEtMp12_qin_b, ScOrEtMp12_qout_d, ScOrEtMp12_qout_e, ScOrEtMp12_qout_v, ScOrEtMp12_qout_b, ScOrEtMp13_qin_d, ScOrEtMp13_qin_e, ScOrEtMp13_qin_v, ScOrEtMp13_qin_b, ScOrEtMp13_qout_d, ScOrEtMp13_qout_e, ScOrEtMp13_qout_v, ScOrEtMp13_qout_b, ScOrEtMp15_qin_d, ScOrEtMp15_qin_e, ScOrEtMp15_qin_v, ScOrEtMp15_qin_b, ScOrEtMp15_qout_d, ScOrEtMp15_qout_e, ScOrEtMp15_qout_v, ScOrEtMp15_qout_b, ScOrEtMp16_qin_d, ScOrEtMp16_qin_e, ScOrEtMp16_qin_v, ScOrEtMp16_qin_b, ScOrEtMp16_qout_d, ScOrEtMp16_qout_e, ScOrEtMp16_qout_v, ScOrEtMp16_qout_b, ScOrEtMp21_qin_d, ScOrEtMp21_qin_e, ScOrEtMp21_qin_v, ScOrEtMp21_qin_b, ScOrEtMp21_qout_d, ScOrEtMp21_qout_e, ScOrEtMp21_qout_v, ScOrEtMp21_qout_b, ScOrEtMp22_qin_d, ScOrEtMp22_qin_e, ScOrEtMp22_qin_v, ScOrEtMp22_qin_b, ScOrEtMp22_qout_d, ScOrEtMp22_qout_e, ScOrEtMp22_qout_v, ScOrEtMp22_qout_b, ScOrEtMp23_qin_d, ScOrEtMp23_qin_e, ScOrEtMp23_qin_v, ScOrEtMp23_qin_b, ScOrEtMp23_qout_d, ScOrEtMp23_qout_e, ScOrEtMp23_qout_v, ScOrEtMp23_qout_b, ScOrEtMp24_qin_d, ScOrEtMp24_qin_e, ScOrEtMp24_qin_v, ScOrEtMp24_qin_b, ScOrEtMp24_qout_d, ScOrEtMp24_qout_e, ScOrEtMp24_qout_v, ScOrEtMp24_qout_b, ScOrEtMp25_qin_d, ScOrEtMp25_qin_e, ScOrEtMp25_qin_v, ScOrEtMp25_qin_b, ScOrEtMp25_qout_d, ScOrEtMp25_qout_e, ScOrEtMp25_qout_v, ScOrEtMp25_qout_b, ScOrEtMp26_qin_d, ScOrEtMp26_qin_e, ScOrEtMp26_qin_v, ScOrEtMp26_qin_b, ScOrEtMp26_qout_d, ScOrEtMp26_qout_e, ScOrEtMp26_qout_v, ScOrEtMp26_qout_b, ScOrEtMp27_qin_d, ScOrEtMp27_qin_e, ScOrEtMp27_qin_v, ScOrEtMp27_qin_b, ScOrEtMp27_qout_d, ScOrEtMp27_qout_e, ScOrEtMp27_qout_v, ScOrEtMp27_qout_b, ScOrEtMp28_qin_d, ScOrEtMp28_qin_e, ScOrEtMp28_qin_v, ScOrEtMp28_qin_b, ScOrEtMp28_qout_d, ScOrEtMp28_qout_e, ScOrEtMp28_qout_v, ScOrEtMp28_qout_b, ScOrEtMp29_qin_d, ScOrEtMp29_qin_e, ScOrEtMp29_qin_v, ScOrEtMp29_qin_b, ScOrEtMp29_qout_d, ScOrEtMp29_qout_e, ScOrEtMp29_qout_v, ScOrEtMp29_qout_b, ScOrEtMp30_qin_d, ScOrEtMp30_qin_e, ScOrEtMp30_qin_v, ScOrEtMp30_qin_b, ScOrEtMp30_qout_d, ScOrEtMp30_qout_e, ScOrEtMp30_qout_v, ScOrEtMp30_qout_b, ScOrEtMp31_qin_d, ScOrEtMp31_qin_e, ScOrEtMp31_qin_v, ScOrEtMp31_qin_b, ScOrEtMp31_qout_d, ScOrEtMp31_qout_e, ScOrEtMp31_qout_v, ScOrEtMp31_qout_b, ScOrEtMp32_qin_d, ScOrEtMp32_qin_e, ScOrEtMp32_qin_v, ScOrEtMp32_qin_b, ScOrEtMp32_qout_d, ScOrEtMp32_qout_e, ScOrEtMp32_qout_v, ScOrEtMp32_qout_b, ScOrEtMp33_qin_d, ScOrEtMp33_qin_e, ScOrEtMp33_qin_v, ScOrEtMp33_qin_b, ScOrEtMp33_qout_d, ScOrEtMp33_qout_e, ScOrEtMp33_qout_v, ScOrEtMp33_qout_b, ScOrEtMp34_qin_d, ScOrEtMp34_qin_e, ScOrEtMp34_qin_v, ScOrEtMp34_qin_b, ScOrEtMp34_qout_d, ScOrEtMp34_qout_e, ScOrEtMp34_qout_v, ScOrEtMp34_qout_b, ScOrEtMp35_qin_d, ScOrEtMp35_qin_e, ScOrEtMp35_qin_v, ScOrEtMp35_qin_b, ScOrEtMp35_qout_d, ScOrEtMp35_qout_e, ScOrEtMp35_qout_v, ScOrEtMp35_qout_b, ScOrEtMp36_qin_d, ScOrEtMp36_qin_e, ScOrEtMp36_qin_v, ScOrEtMp36_qin_b, ScOrEtMp36_qout_d, ScOrEtMp36_qout_e, ScOrEtMp36_qout_v, ScOrEtMp36_qout_b, ScOrEtMp37_qin_d, ScOrEtMp37_qin_e, ScOrEtMp37_qin_v, ScOrEtMp37_qin_b, ScOrEtMp37_qout_d, ScOrEtMp37_qout_e, ScOrEtMp37_qout_v, ScOrEtMp37_qout_b, ScOrEtMp38_qin_d, ScOrEtMp38_qin_e, ScOrEtMp38_qin_v, ScOrEtMp38_qin_b, ScOrEtMp38_qout_d, ScOrEtMp38_qout_e, ScOrEtMp38_qout_v, ScOrEtMp38_qout_b, ScOrEtMp39_qin_d, ScOrEtMp39_qin_e, ScOrEtMp39_qin_v, ScOrEtMp39_qin_b, ScOrEtMp39_qout_d, ScOrEtMp39_qout_e, ScOrEtMp39_qout_v, ScOrEtMp39_qout_b, ScOrEtMp40_qin_d, ScOrEtMp40_qin_e, ScOrEtMp40_qin_v, ScOrEtMp40_qin_b, ScOrEtMp40_qout_d, ScOrEtMp40_qout_e, ScOrEtMp40_qout_v, ScOrEtMp40_qout_b, ScOrEtMp41_qin_d, ScOrEtMp41_qin_e, ScOrEtMp41_qin_v, ScOrEtMp41_qin_b, ScOrEtMp41_qout_d, ScOrEtMp41_qout_e, ScOrEtMp41_qout_v, ScOrEtMp41_qout_b, ScOrEtMp42_qin_d, ScOrEtMp42_qin_e, ScOrEtMp42_qin_v, ScOrEtMp42_qin_b, ScOrEtMp42_qout_d, ScOrEtMp42_qout_e, ScOrEtMp42_qout_v, ScOrEtMp42_qout_b, ScOrEtMp43_qin_d, ScOrEtMp43_qin_e, ScOrEtMp43_qin_v, ScOrEtMp43_qin_b, ScOrEtMp43_qout_d, ScOrEtMp43_qout_e, ScOrEtMp43_qout_v, ScOrEtMp43_qout_b, ScOrEtMp44_qin_d, ScOrEtMp44_qin_e, ScOrEtMp44_qin_v, ScOrEtMp44_qin_b, ScOrEtMp44_qout_d, ScOrEtMp44_qout_e, ScOrEtMp44_qout_v, ScOrEtMp44_qout_b, ScOrEtMp55_qin_d, ScOrEtMp55_qin_e, ScOrEtMp55_qin_v, ScOrEtMp55_qin_b, ScOrEtMp55_qout_d, ScOrEtMp55_qout_e, ScOrEtMp55_qout_v, ScOrEtMp55_qout_b, ScOrEtMp56_qin_d, ScOrEtMp56_qin_e, ScOrEtMp56_qin_v, ScOrEtMp56_qin_b, ScOrEtMp56_qout_d, ScOrEtMp56_qout_e, ScOrEtMp56_qout_v, ScOrEtMp56_qout_b);

  input  clock;
  input  reset;

  input  [8:0] outA_qin_d;
  input  outA_qin_e;
  input  outA_qin_v;
  output outA_qin_b;
  output [8:0] outA_qout_d;
  output outA_qout_e;
  output outA_qout_v;
  input  outA_qout_b;
  input  [8:0] outB_qin_d;
  input  outB_qin_e;
  input  outB_qin_v;
  output outB_qin_b;
  output [8:0] outB_qout_d;
  output outB_qout_e;
  output outB_qout_v;
  input  outB_qout_b;
  input  [8:0] outC_qin_d;
  input  outC_qin_e;
  input  outC_qin_v;
  output outC_qin_b;
  output [8:0] outC_qout_d;
  output outC_qout_e;
  output outC_qout_v;
  input  outC_qout_b;
  input  [8:0] outD_qin_d;
  input  outD_qin_e;
  input  outD_qin_v;
  output outD_qin_b;
  output [8:0] outD_qout_d;
  output outD_qout_e;
  output outD_qout_v;
  input  outD_qout_b;
  input  [8:0] outE_qin_d;
  input  outE_qin_e;
  input  outE_qin_v;
  output outE_qin_b;
  output [8:0] outE_qout_d;
  output outE_qout_e;
  output outE_qout_v;
  input  outE_qout_b;
  input  [8:0] outF_qin_d;
  input  outF_qin_e;
  input  outF_qin_v;
  output outF_qin_b;
  output [8:0] outF_qout_d;
  output outF_qout_e;
  output outF_qout_v;
  input  outF_qout_b;
  input  [8:0] outG_qin_d;
  input  outG_qin_e;
  input  outG_qin_v;
  output outG_qin_b;
  output [8:0] outG_qout_d;
  output outG_qout_e;
  output outG_qout_v;
  input  outG_qout_b;
  input  [8:0] outH_qin_d;
  input  outH_qin_e;
  input  outH_qin_v;
  output outH_qin_b;
  output [8:0] outH_qout_d;
  output outH_qout_e;
  output outH_qout_v;
  input  outH_qout_b;
  input  [15:0] ScOrEtMp1_qin_d;
  input  ScOrEtMp1_qin_e;
  input  ScOrEtMp1_qin_v;
  output ScOrEtMp1_qin_b;
  output [15:0] ScOrEtMp1_qout_d;
  output ScOrEtMp1_qout_e;
  output ScOrEtMp1_qout_v;
  input  ScOrEtMp1_qout_b;
  input  [15:0] ScOrEtMp2_qin_d;
  input  ScOrEtMp2_qin_e;
  input  ScOrEtMp2_qin_v;
  output ScOrEtMp2_qin_b;
  output [15:0] ScOrEtMp2_qout_d;
  output ScOrEtMp2_qout_e;
  output ScOrEtMp2_qout_v;
  input  ScOrEtMp2_qout_b;
  input  [15:0] ScOrEtMp3_qin_d;
  input  ScOrEtMp3_qin_e;
  input  ScOrEtMp3_qin_v;
  output ScOrEtMp3_qin_b;
  output [15:0] ScOrEtMp3_qout_d;
  output ScOrEtMp3_qout_e;
  output ScOrEtMp3_qout_v;
  input  ScOrEtMp3_qout_b;
  input  [15:0] ScOrEtMp4_qin_d;
  input  ScOrEtMp4_qin_e;
  input  ScOrEtMp4_qin_v;
  output ScOrEtMp4_qin_b;
  output [15:0] ScOrEtMp4_qout_d;
  output ScOrEtMp4_qout_e;
  output ScOrEtMp4_qout_v;
  input  ScOrEtMp4_qout_b;
  input  [15:0] ScOrEtMp5_qin_d;
  input  ScOrEtMp5_qin_e;
  input  ScOrEtMp5_qin_v;
  output ScOrEtMp5_qin_b;
  output [15:0] ScOrEtMp5_qout_d;
  output ScOrEtMp5_qout_e;
  output ScOrEtMp5_qout_v;
  input  ScOrEtMp5_qout_b;
  input  [15:0] ScOrEtMp6_qin_d;
  input  ScOrEtMp6_qin_e;
  input  ScOrEtMp6_qin_v;
  output ScOrEtMp6_qin_b;
  output [15:0] ScOrEtMp6_qout_d;
  output ScOrEtMp6_qout_e;
  output ScOrEtMp6_qout_v;
  input  ScOrEtMp6_qout_b;
  input  [15:0] ScOrEtMp7_qin_d;
  input  ScOrEtMp7_qin_e;
  input  ScOrEtMp7_qin_v;
  output ScOrEtMp7_qin_b;
  output [15:0] ScOrEtMp7_qout_d;
  output ScOrEtMp7_qout_e;
  output ScOrEtMp7_qout_v;
  input  ScOrEtMp7_qout_b;
  input  [15:0] ScOrEtMp8_qin_d;
  input  ScOrEtMp8_qin_e;
  input  ScOrEtMp8_qin_v;
  output ScOrEtMp8_qin_b;
  output [15:0] ScOrEtMp8_qout_d;
  output ScOrEtMp8_qout_e;
  output ScOrEtMp8_qout_v;
  input  ScOrEtMp8_qout_b;
  input  [15:0] ScOrEtMp9_qin_d;
  input  ScOrEtMp9_qin_e;
  input  ScOrEtMp9_qin_v;
  output ScOrEtMp9_qin_b;
  output [15:0] ScOrEtMp9_qout_d;
  output ScOrEtMp9_qout_e;
  output ScOrEtMp9_qout_v;
  input  ScOrEtMp9_qout_b;
  input  [15:0] ScOrEtMp10_qin_d;
  input  ScOrEtMp10_qin_e;
  input  ScOrEtMp10_qin_v;
  output ScOrEtMp10_qin_b;
  output [15:0] ScOrEtMp10_qout_d;
  output ScOrEtMp10_qout_e;
  output ScOrEtMp10_qout_v;
  input  ScOrEtMp10_qout_b;
  input  [15:0] ScOrEtMp11_qin_d;
  input  ScOrEtMp11_qin_e;
  input  ScOrEtMp11_qin_v;
  output ScOrEtMp11_qin_b;
  output [15:0] ScOrEtMp11_qout_d;
  output ScOrEtMp11_qout_e;
  output ScOrEtMp11_qout_v;
  input  ScOrEtMp11_qout_b;
  input  [7:0] ScOrEtMp12_qin_d;
  input  ScOrEtMp12_qin_e;
  input  ScOrEtMp12_qin_v;
  output ScOrEtMp12_qin_b;
  output [7:0] ScOrEtMp12_qout_d;
  output ScOrEtMp12_qout_e;
  output ScOrEtMp12_qout_v;
  input  ScOrEtMp12_qout_b;
  input  [7:0] ScOrEtMp13_qin_d;
  input  ScOrEtMp13_qin_e;
  input  ScOrEtMp13_qin_v;
  output ScOrEtMp13_qin_b;
  output [7:0] ScOrEtMp13_qout_d;
  output ScOrEtMp13_qout_e;
  output ScOrEtMp13_qout_v;
  input  ScOrEtMp13_qout_b;
  input  [7:0] ScOrEtMp15_qin_d;
  input  ScOrEtMp15_qin_e;
  input  ScOrEtMp15_qin_v;
  output ScOrEtMp15_qin_b;
  output [7:0] ScOrEtMp15_qout_d;
  output ScOrEtMp15_qout_e;
  output ScOrEtMp15_qout_v;
  input  ScOrEtMp15_qout_b;
  input  [7:0] ScOrEtMp16_qin_d;
  input  ScOrEtMp16_qin_e;
  input  ScOrEtMp16_qin_v;
  output ScOrEtMp16_qin_b;
  output [7:0] ScOrEtMp16_qout_d;
  output ScOrEtMp16_qout_e;
  output ScOrEtMp16_qout_v;
  input  ScOrEtMp16_qout_b;
  input  [15:0] ScOrEtMp21_qin_d;
  input  ScOrEtMp21_qin_e;
  input  ScOrEtMp21_qin_v;
  output ScOrEtMp21_qin_b;
  output [15:0] ScOrEtMp21_qout_d;
  output ScOrEtMp21_qout_e;
  output ScOrEtMp21_qout_v;
  input  ScOrEtMp21_qout_b;
  input  [15:0] ScOrEtMp22_qin_d;
  input  ScOrEtMp22_qin_e;
  input  ScOrEtMp22_qin_v;
  output ScOrEtMp22_qin_b;
  output [15:0] ScOrEtMp22_qout_d;
  output ScOrEtMp22_qout_e;
  output ScOrEtMp22_qout_v;
  input  ScOrEtMp22_qout_b;
  input  [15:0] ScOrEtMp23_qin_d;
  input  ScOrEtMp23_qin_e;
  input  ScOrEtMp23_qin_v;
  output ScOrEtMp23_qin_b;
  output [15:0] ScOrEtMp23_qout_d;
  output ScOrEtMp23_qout_e;
  output ScOrEtMp23_qout_v;
  input  ScOrEtMp23_qout_b;
  input  [15:0] ScOrEtMp24_qin_d;
  input  ScOrEtMp24_qin_e;
  input  ScOrEtMp24_qin_v;
  output ScOrEtMp24_qin_b;
  output [15:0] ScOrEtMp24_qout_d;
  output ScOrEtMp24_qout_e;
  output ScOrEtMp24_qout_v;
  input  ScOrEtMp24_qout_b;
  input  [15:0] ScOrEtMp25_qin_d;
  input  ScOrEtMp25_qin_e;
  input  ScOrEtMp25_qin_v;
  output ScOrEtMp25_qin_b;
  output [15:0] ScOrEtMp25_qout_d;
  output ScOrEtMp25_qout_e;
  output ScOrEtMp25_qout_v;
  input  ScOrEtMp25_qout_b;
  input  [15:0] ScOrEtMp26_qin_d;
  input  ScOrEtMp26_qin_e;
  input  ScOrEtMp26_qin_v;
  output ScOrEtMp26_qin_b;
  output [15:0] ScOrEtMp26_qout_d;
  output ScOrEtMp26_qout_e;
  output ScOrEtMp26_qout_v;
  input  ScOrEtMp26_qout_b;
  input  [15:0] ScOrEtMp27_qin_d;
  input  ScOrEtMp27_qin_e;
  input  ScOrEtMp27_qin_v;
  output ScOrEtMp27_qin_b;
  output [15:0] ScOrEtMp27_qout_d;
  output ScOrEtMp27_qout_e;
  output ScOrEtMp27_qout_v;
  input  ScOrEtMp27_qout_b;
  input  [15:0] ScOrEtMp28_qin_d;
  input  ScOrEtMp28_qin_e;
  input  ScOrEtMp28_qin_v;
  output ScOrEtMp28_qin_b;
  output [15:0] ScOrEtMp28_qout_d;
  output ScOrEtMp28_qout_e;
  output ScOrEtMp28_qout_v;
  input  ScOrEtMp28_qout_b;
  input  [15:0] ScOrEtMp29_qin_d;
  input  ScOrEtMp29_qin_e;
  input  ScOrEtMp29_qin_v;
  output ScOrEtMp29_qin_b;
  output [15:0] ScOrEtMp29_qout_d;
  output ScOrEtMp29_qout_e;
  output ScOrEtMp29_qout_v;
  input  ScOrEtMp29_qout_b;
  input  [15:0] ScOrEtMp30_qin_d;
  input  ScOrEtMp30_qin_e;
  input  ScOrEtMp30_qin_v;
  output ScOrEtMp30_qin_b;
  output [15:0] ScOrEtMp30_qout_d;
  output ScOrEtMp30_qout_e;
  output ScOrEtMp30_qout_v;
  input  ScOrEtMp30_qout_b;
  input  [15:0] ScOrEtMp31_qin_d;
  input  ScOrEtMp31_qin_e;
  input  ScOrEtMp31_qin_v;
  output ScOrEtMp31_qin_b;
  output [15:0] ScOrEtMp31_qout_d;
  output ScOrEtMp31_qout_e;
  output ScOrEtMp31_qout_v;
  input  ScOrEtMp31_qout_b;
  input  [15:0] ScOrEtMp32_qin_d;
  input  ScOrEtMp32_qin_e;
  input  ScOrEtMp32_qin_v;
  output ScOrEtMp32_qin_b;
  output [15:0] ScOrEtMp32_qout_d;
  output ScOrEtMp32_qout_e;
  output ScOrEtMp32_qout_v;
  input  ScOrEtMp32_qout_b;
  input  [15:0] ScOrEtMp33_qin_d;
  input  ScOrEtMp33_qin_e;
  input  ScOrEtMp33_qin_v;
  output ScOrEtMp33_qin_b;
  output [15:0] ScOrEtMp33_qout_d;
  output ScOrEtMp33_qout_e;
  output ScOrEtMp33_qout_v;
  input  ScOrEtMp33_qout_b;
  input  [15:0] ScOrEtMp34_qin_d;
  input  ScOrEtMp34_qin_e;
  input  ScOrEtMp34_qin_v;
  output ScOrEtMp34_qin_b;
  output [15:0] ScOrEtMp34_qout_d;
  output ScOrEtMp34_qout_e;
  output ScOrEtMp34_qout_v;
  input  ScOrEtMp34_qout_b;
  input  [15:0] ScOrEtMp35_qin_d;
  input  ScOrEtMp35_qin_e;
  input  ScOrEtMp35_qin_v;
  output ScOrEtMp35_qin_b;
  output [15:0] ScOrEtMp35_qout_d;
  output ScOrEtMp35_qout_e;
  output ScOrEtMp35_qout_v;
  input  ScOrEtMp35_qout_b;
  input  [15:0] ScOrEtMp36_qin_d;
  input  ScOrEtMp36_qin_e;
  input  ScOrEtMp36_qin_v;
  output ScOrEtMp36_qin_b;
  output [15:0] ScOrEtMp36_qout_d;
  output ScOrEtMp36_qout_e;
  output ScOrEtMp36_qout_v;
  input  ScOrEtMp36_qout_b;
  input  [8:0] ScOrEtMp37_qin_d;
  input  ScOrEtMp37_qin_e;
  input  ScOrEtMp37_qin_v;
  output ScOrEtMp37_qin_b;
  output [8:0] ScOrEtMp37_qout_d;
  output ScOrEtMp37_qout_e;
  output ScOrEtMp37_qout_v;
  input  ScOrEtMp37_qout_b;
  input  [8:0] ScOrEtMp38_qin_d;
  input  ScOrEtMp38_qin_e;
  input  ScOrEtMp38_qin_v;
  output ScOrEtMp38_qin_b;
  output [8:0] ScOrEtMp38_qout_d;
  output ScOrEtMp38_qout_e;
  output ScOrEtMp38_qout_v;
  input  ScOrEtMp38_qout_b;
  input  [8:0] ScOrEtMp39_qin_d;
  input  ScOrEtMp39_qin_e;
  input  ScOrEtMp39_qin_v;
  output ScOrEtMp39_qin_b;
  output [8:0] ScOrEtMp39_qout_d;
  output ScOrEtMp39_qout_e;
  output ScOrEtMp39_qout_v;
  input  ScOrEtMp39_qout_b;
  input  [8:0] ScOrEtMp40_qin_d;
  input  ScOrEtMp40_qin_e;
  input  ScOrEtMp40_qin_v;
  output ScOrEtMp40_qin_b;
  output [8:0] ScOrEtMp40_qout_d;
  output ScOrEtMp40_qout_e;
  output ScOrEtMp40_qout_v;
  input  ScOrEtMp40_qout_b;
  input  [8:0] ScOrEtMp41_qin_d;
  input  ScOrEtMp41_qin_e;
  input  ScOrEtMp41_qin_v;
  output ScOrEtMp41_qin_b;
  output [8:0] ScOrEtMp41_qout_d;
  output ScOrEtMp41_qout_e;
  output ScOrEtMp41_qout_v;
  input  ScOrEtMp41_qout_b;
  input  [8:0] ScOrEtMp42_qin_d;
  input  ScOrEtMp42_qin_e;
  input  ScOrEtMp42_qin_v;
  output ScOrEtMp42_qin_b;
  output [8:0] ScOrEtMp42_qout_d;
  output ScOrEtMp42_qout_e;
  output ScOrEtMp42_qout_v;
  input  ScOrEtMp42_qout_b;
  input  [8:0] ScOrEtMp43_qin_d;
  input  ScOrEtMp43_qin_e;
  input  ScOrEtMp43_qin_v;
  output ScOrEtMp43_qin_b;
  output [8:0] ScOrEtMp43_qout_d;
  output ScOrEtMp43_qout_e;
  output ScOrEtMp43_qout_v;
  input  ScOrEtMp43_qout_b;
  input  [8:0] ScOrEtMp44_qin_d;
  input  ScOrEtMp44_qin_e;
  input  ScOrEtMp44_qin_v;
  output ScOrEtMp44_qin_b;
  output [8:0] ScOrEtMp44_qout_d;
  output ScOrEtMp44_qout_e;
  output ScOrEtMp44_qout_v;
  input  ScOrEtMp44_qout_b;
  input  [31:0] ScOrEtMp55_qin_d;
  input  ScOrEtMp55_qin_e;
  input  ScOrEtMp55_qin_v;
  output ScOrEtMp55_qin_b;
  output [31:0] ScOrEtMp55_qout_d;
  output ScOrEtMp55_qout_e;
  output ScOrEtMp55_qout_v;
  input  ScOrEtMp55_qout_b;
  input  [63:0] ScOrEtMp56_qin_d;
  input  ScOrEtMp56_qin_e;
  input  ScOrEtMp56_qin_v;
  output ScOrEtMp56_qin_b;
  output [63:0] ScOrEtMp56_qout_d;
  output ScOrEtMp56_qout_e;
  output ScOrEtMp56_qout_v;
  input  ScOrEtMp56_qout_b;

  Q_wire #(0, 10) q_outA (clock, reset, {outA_qin_d, outA_qin_e}, outA_qin_v, outA_qin_b, {outA_qout_d, outA_qout_e}, outA_qout_v, outA_qout_b);
  Q_wire #(0, 10) q_outB (clock, reset, {outB_qin_d, outB_qin_e}, outB_qin_v, outB_qin_b, {outB_qout_d, outB_qout_e}, outB_qout_v, outB_qout_b);
  Q_wire #(0, 10) q_outC (clock, reset, {outC_qin_d, outC_qin_e}, outC_qin_v, outC_qin_b, {outC_qout_d, outC_qout_e}, outC_qout_v, outC_qout_b);
  Q_wire #(0, 10) q_outD (clock, reset, {outD_qin_d, outD_qin_e}, outD_qin_v, outD_qin_b, {outD_qout_d, outD_qout_e}, outD_qout_v, outD_qout_b);
  Q_wire #(0, 10) q_outE (clock, reset, {outE_qin_d, outE_qin_e}, outE_qin_v, outE_qin_b, {outE_qout_d, outE_qout_e}, outE_qout_v, outE_qout_b);
  Q_wire #(0, 10) q_outF (clock, reset, {outF_qin_d, outF_qin_e}, outF_qin_v, outF_qin_b, {outF_qout_d, outF_qout_e}, outF_qout_v, outF_qout_b);
  Q_wire #(0, 10) q_outG (clock, reset, {outG_qin_d, outG_qin_e}, outG_qin_v, outG_qin_b, {outG_qout_d, outG_qout_e}, outG_qout_v, outG_qout_b);
  Q_wire #(0, 10) q_outH (clock, reset, {outH_qin_d, outH_qin_e}, outH_qin_v, outH_qin_b, {outH_qout_d, outH_qout_e}, outH_qout_v, outH_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp1 (clock, reset, {ScOrEtMp1_qin_d, ScOrEtMp1_qin_e}, ScOrEtMp1_qin_v, ScOrEtMp1_qin_b, {ScOrEtMp1_qout_d, ScOrEtMp1_qout_e}, ScOrEtMp1_qout_v, ScOrEtMp1_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp2 (clock, reset, {ScOrEtMp2_qin_d, ScOrEtMp2_qin_e}, ScOrEtMp2_qin_v, ScOrEtMp2_qin_b, {ScOrEtMp2_qout_d, ScOrEtMp2_qout_e}, ScOrEtMp2_qout_v, ScOrEtMp2_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp3 (clock, reset, {ScOrEtMp3_qin_d, ScOrEtMp3_qin_e}, ScOrEtMp3_qin_v, ScOrEtMp3_qin_b, {ScOrEtMp3_qout_d, ScOrEtMp3_qout_e}, ScOrEtMp3_qout_v, ScOrEtMp3_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp4 (clock, reset, {ScOrEtMp4_qin_d, ScOrEtMp4_qin_e}, ScOrEtMp4_qin_v, ScOrEtMp4_qin_b, {ScOrEtMp4_qout_d, ScOrEtMp4_qout_e}, ScOrEtMp4_qout_v, ScOrEtMp4_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp5 (clock, reset, {ScOrEtMp5_qin_d, ScOrEtMp5_qin_e}, ScOrEtMp5_qin_v, ScOrEtMp5_qin_b, {ScOrEtMp5_qout_d, ScOrEtMp5_qout_e}, ScOrEtMp5_qout_v, ScOrEtMp5_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp6 (clock, reset, {ScOrEtMp6_qin_d, ScOrEtMp6_qin_e}, ScOrEtMp6_qin_v, ScOrEtMp6_qin_b, {ScOrEtMp6_qout_d, ScOrEtMp6_qout_e}, ScOrEtMp6_qout_v, ScOrEtMp6_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp7 (clock, reset, {ScOrEtMp7_qin_d, ScOrEtMp7_qin_e}, ScOrEtMp7_qin_v, ScOrEtMp7_qin_b, {ScOrEtMp7_qout_d, ScOrEtMp7_qout_e}, ScOrEtMp7_qout_v, ScOrEtMp7_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp8 (clock, reset, {ScOrEtMp8_qin_d, ScOrEtMp8_qin_e}, ScOrEtMp8_qin_v, ScOrEtMp8_qin_b, {ScOrEtMp8_qout_d, ScOrEtMp8_qout_e}, ScOrEtMp8_qout_v, ScOrEtMp8_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp9 (clock, reset, {ScOrEtMp9_qin_d, ScOrEtMp9_qin_e}, ScOrEtMp9_qin_v, ScOrEtMp9_qin_b, {ScOrEtMp9_qout_d, ScOrEtMp9_qout_e}, ScOrEtMp9_qout_v, ScOrEtMp9_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp10 (clock, reset, {ScOrEtMp10_qin_d, ScOrEtMp10_qin_e}, ScOrEtMp10_qin_v, ScOrEtMp10_qin_b, {ScOrEtMp10_qout_d, ScOrEtMp10_qout_e}, ScOrEtMp10_qout_v, ScOrEtMp10_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp11 (clock, reset, {ScOrEtMp11_qin_d, ScOrEtMp11_qin_e}, ScOrEtMp11_qin_v, ScOrEtMp11_qin_b, {ScOrEtMp11_qout_d, ScOrEtMp11_qout_e}, ScOrEtMp11_qout_v, ScOrEtMp11_qout_b);
  Q_wire #(0, 9) q_ScOrEtMp12 (clock, reset, {ScOrEtMp12_qin_d, ScOrEtMp12_qin_e}, ScOrEtMp12_qin_v, ScOrEtMp12_qin_b, {ScOrEtMp12_qout_d, ScOrEtMp12_qout_e}, ScOrEtMp12_qout_v, ScOrEtMp12_qout_b);
  Q_wire #(0, 9) q_ScOrEtMp13 (clock, reset, {ScOrEtMp13_qin_d, ScOrEtMp13_qin_e}, ScOrEtMp13_qin_v, ScOrEtMp13_qin_b, {ScOrEtMp13_qout_d, ScOrEtMp13_qout_e}, ScOrEtMp13_qout_v, ScOrEtMp13_qout_b);
  Q_wire #(0, 9) q_ScOrEtMp15 (clock, reset, {ScOrEtMp15_qin_d, ScOrEtMp15_qin_e}, ScOrEtMp15_qin_v, ScOrEtMp15_qin_b, {ScOrEtMp15_qout_d, ScOrEtMp15_qout_e}, ScOrEtMp15_qout_v, ScOrEtMp15_qout_b);
  Q_wire #(0, 9) q_ScOrEtMp16 (clock, reset, {ScOrEtMp16_qin_d, ScOrEtMp16_qin_e}, ScOrEtMp16_qin_v, ScOrEtMp16_qin_b, {ScOrEtMp16_qout_d, ScOrEtMp16_qout_e}, ScOrEtMp16_qout_v, ScOrEtMp16_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp21 (clock, reset, {ScOrEtMp21_qin_d, ScOrEtMp21_qin_e}, ScOrEtMp21_qin_v, ScOrEtMp21_qin_b, {ScOrEtMp21_qout_d, ScOrEtMp21_qout_e}, ScOrEtMp21_qout_v, ScOrEtMp21_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp22 (clock, reset, {ScOrEtMp22_qin_d, ScOrEtMp22_qin_e}, ScOrEtMp22_qin_v, ScOrEtMp22_qin_b, {ScOrEtMp22_qout_d, ScOrEtMp22_qout_e}, ScOrEtMp22_qout_v, ScOrEtMp22_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp23 (clock, reset, {ScOrEtMp23_qin_d, ScOrEtMp23_qin_e}, ScOrEtMp23_qin_v, ScOrEtMp23_qin_b, {ScOrEtMp23_qout_d, ScOrEtMp23_qout_e}, ScOrEtMp23_qout_v, ScOrEtMp23_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp24 (clock, reset, {ScOrEtMp24_qin_d, ScOrEtMp24_qin_e}, ScOrEtMp24_qin_v, ScOrEtMp24_qin_b, {ScOrEtMp24_qout_d, ScOrEtMp24_qout_e}, ScOrEtMp24_qout_v, ScOrEtMp24_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp25 (clock, reset, {ScOrEtMp25_qin_d, ScOrEtMp25_qin_e}, ScOrEtMp25_qin_v, ScOrEtMp25_qin_b, {ScOrEtMp25_qout_d, ScOrEtMp25_qout_e}, ScOrEtMp25_qout_v, ScOrEtMp25_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp26 (clock, reset, {ScOrEtMp26_qin_d, ScOrEtMp26_qin_e}, ScOrEtMp26_qin_v, ScOrEtMp26_qin_b, {ScOrEtMp26_qout_d, ScOrEtMp26_qout_e}, ScOrEtMp26_qout_v, ScOrEtMp26_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp27 (clock, reset, {ScOrEtMp27_qin_d, ScOrEtMp27_qin_e}, ScOrEtMp27_qin_v, ScOrEtMp27_qin_b, {ScOrEtMp27_qout_d, ScOrEtMp27_qout_e}, ScOrEtMp27_qout_v, ScOrEtMp27_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp28 (clock, reset, {ScOrEtMp28_qin_d, ScOrEtMp28_qin_e}, ScOrEtMp28_qin_v, ScOrEtMp28_qin_b, {ScOrEtMp28_qout_d, ScOrEtMp28_qout_e}, ScOrEtMp28_qout_v, ScOrEtMp28_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp29 (clock, reset, {ScOrEtMp29_qin_d, ScOrEtMp29_qin_e}, ScOrEtMp29_qin_v, ScOrEtMp29_qin_b, {ScOrEtMp29_qout_d, ScOrEtMp29_qout_e}, ScOrEtMp29_qout_v, ScOrEtMp29_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp30 (clock, reset, {ScOrEtMp30_qin_d, ScOrEtMp30_qin_e}, ScOrEtMp30_qin_v, ScOrEtMp30_qin_b, {ScOrEtMp30_qout_d, ScOrEtMp30_qout_e}, ScOrEtMp30_qout_v, ScOrEtMp30_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp31 (clock, reset, {ScOrEtMp31_qin_d, ScOrEtMp31_qin_e}, ScOrEtMp31_qin_v, ScOrEtMp31_qin_b, {ScOrEtMp31_qout_d, ScOrEtMp31_qout_e}, ScOrEtMp31_qout_v, ScOrEtMp31_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp32 (clock, reset, {ScOrEtMp32_qin_d, ScOrEtMp32_qin_e}, ScOrEtMp32_qin_v, ScOrEtMp32_qin_b, {ScOrEtMp32_qout_d, ScOrEtMp32_qout_e}, ScOrEtMp32_qout_v, ScOrEtMp32_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp33 (clock, reset, {ScOrEtMp33_qin_d, ScOrEtMp33_qin_e}, ScOrEtMp33_qin_v, ScOrEtMp33_qin_b, {ScOrEtMp33_qout_d, ScOrEtMp33_qout_e}, ScOrEtMp33_qout_v, ScOrEtMp33_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp34 (clock, reset, {ScOrEtMp34_qin_d, ScOrEtMp34_qin_e}, ScOrEtMp34_qin_v, ScOrEtMp34_qin_b, {ScOrEtMp34_qout_d, ScOrEtMp34_qout_e}, ScOrEtMp34_qout_v, ScOrEtMp34_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp35 (clock, reset, {ScOrEtMp35_qin_d, ScOrEtMp35_qin_e}, ScOrEtMp35_qin_v, ScOrEtMp35_qin_b, {ScOrEtMp35_qout_d, ScOrEtMp35_qout_e}, ScOrEtMp35_qout_v, ScOrEtMp35_qout_b);
  Q_wire #(0, 17) q_ScOrEtMp36 (clock, reset, {ScOrEtMp36_qin_d, ScOrEtMp36_qin_e}, ScOrEtMp36_qin_v, ScOrEtMp36_qin_b, {ScOrEtMp36_qout_d, ScOrEtMp36_qout_e}, ScOrEtMp36_qout_v, ScOrEtMp36_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp37 (clock, reset, {ScOrEtMp37_qin_d, ScOrEtMp37_qin_e}, ScOrEtMp37_qin_v, ScOrEtMp37_qin_b, {ScOrEtMp37_qout_d, ScOrEtMp37_qout_e}, ScOrEtMp37_qout_v, ScOrEtMp37_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp38 (clock, reset, {ScOrEtMp38_qin_d, ScOrEtMp38_qin_e}, ScOrEtMp38_qin_v, ScOrEtMp38_qin_b, {ScOrEtMp38_qout_d, ScOrEtMp38_qout_e}, ScOrEtMp38_qout_v, ScOrEtMp38_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp39 (clock, reset, {ScOrEtMp39_qin_d, ScOrEtMp39_qin_e}, ScOrEtMp39_qin_v, ScOrEtMp39_qin_b, {ScOrEtMp39_qout_d, ScOrEtMp39_qout_e}, ScOrEtMp39_qout_v, ScOrEtMp39_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp40 (clock, reset, {ScOrEtMp40_qin_d, ScOrEtMp40_qin_e}, ScOrEtMp40_qin_v, ScOrEtMp40_qin_b, {ScOrEtMp40_qout_d, ScOrEtMp40_qout_e}, ScOrEtMp40_qout_v, ScOrEtMp40_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp41 (clock, reset, {ScOrEtMp41_qin_d, ScOrEtMp41_qin_e}, ScOrEtMp41_qin_v, ScOrEtMp41_qin_b, {ScOrEtMp41_qout_d, ScOrEtMp41_qout_e}, ScOrEtMp41_qout_v, ScOrEtMp41_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp42 (clock, reset, {ScOrEtMp42_qin_d, ScOrEtMp42_qin_e}, ScOrEtMp42_qin_v, ScOrEtMp42_qin_b, {ScOrEtMp42_qout_d, ScOrEtMp42_qout_e}, ScOrEtMp42_qout_v, ScOrEtMp42_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp43 (clock, reset, {ScOrEtMp43_qin_d, ScOrEtMp43_qin_e}, ScOrEtMp43_qin_v, ScOrEtMp43_qin_b, {ScOrEtMp43_qout_d, ScOrEtMp43_qout_e}, ScOrEtMp43_qout_v, ScOrEtMp43_qout_b);
  Q_wire #(0, 10) q_ScOrEtMp44 (clock, reset, {ScOrEtMp44_qin_d, ScOrEtMp44_qin_e}, ScOrEtMp44_qin_v, ScOrEtMp44_qin_b, {ScOrEtMp44_qout_d, ScOrEtMp44_qout_e}, ScOrEtMp44_qout_v, ScOrEtMp44_qout_b);
  Q_wire #(0, 33) q_ScOrEtMp55 (clock, reset, {ScOrEtMp55_qin_d, ScOrEtMp55_qin_e}, ScOrEtMp55_qin_v, ScOrEtMp55_qin_b, {ScOrEtMp55_qout_d, ScOrEtMp55_qout_e}, ScOrEtMp55_qout_v, ScOrEtMp55_qout_b);
  Q_wire #(0, 65) q_ScOrEtMp56 (clock, reset, {ScOrEtMp56_qin_d, ScOrEtMp56_qin_e}, ScOrEtMp56_qin_v, ScOrEtMp56_qin_b, {ScOrEtMp56_qout_d, ScOrEtMp56_qout_e}, ScOrEtMp56_qout_v, ScOrEtMp56_qout_b);

endmodule  // JPEG_dec_d1_ScOrEtMp0_q
