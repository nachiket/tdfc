// Verilog page module without input queues or fsms for _page_illm_d1_ScOrEtMp48
// Emitted by ../../../tdfc version 1.160, Mon Aug 24 17:52:43 2009

`include "_page_illm_d1_ScOrEtMp48_q.v"
`include "illm_d1_ScOrEtMp48_dp.v"

module illm_d1_ScOrEtMp48_fsm (clock, reset, a0_e, a0_v, a0_b, a1_e, a1_v, a1_b, a2_e, a2_v, a2_b, a3_e, a3_v, a3_b, a4_e, a4_v, a4_b, a5_e, a5_v, a5_b, a6_e, a6_v, a6_b, a7_e, a7_v, a7_b, b0_e, b0_v, b0_b, b1_e, b1_v, b1_b, b2_e, b2_v, b2_b, b3_e, b3_v, b3_b, b4_e, b4_v, b4_b, b5_e, b5_v, b5_b, b6_e, b6_v, b6_b, b7_e, b7_v, b7_b, statecase) /* synthesis syn_black_box */ ;

  input  clock;
  input  reset;

  input  a0_e;
  input  a0_v;
  output a0_b;
  input  a1_e;
  input  a1_v;
  output a1_b;
  input  a2_e;
  input  a2_v;
  output a2_b;
  input  a3_e;
  input  a3_v;
  output a3_b;
  input  a4_e;
  input  a4_v;
  output a4_b;
  input  a5_e;
  input  a5_v;
  output a5_b;
  input  a6_e;
  input  a6_v;
  output a6_b;
  input  a7_e;
  input  a7_v;
  output a7_b;
  output b0_e;
  output b0_v;
  input  b0_b;
  output b1_e;
  output b1_v;
  input  b1_b;
  output b2_e;
  output b2_v;
  input  b2_b;
  output b3_e;
  output b3_v;
  input  b3_b;
  output b4_e;
  output b4_v;
  input  b4_b;
  output b5_e;
  output b5_v;
  input  b5_b;
  output b6_e;
  output b6_v;
  input  b6_b;
  output b7_e;
  output b7_v;
  input  b7_b;

  output statecase;

endmodule  // illm_d1_ScOrEtMp48_fsm

module illm_d1_ScOrEtMp48 (clock, reset, a0_d, a0_e, a0_v, a0_b, a1_d, a1_e, a1_v, a1_b, a2_d, a2_e, a2_v, a2_b, a3_d, a3_e, a3_v, a3_b, a4_d, a4_e, a4_v, a4_b, a5_d, a5_e, a5_v, a5_b, a6_d, a6_e, a6_v, a6_b, a7_d, a7_e, a7_v, a7_b, b0_d, b0_e, b0_v, b0_b, b1_d, b1_e, b1_v, b1_b, b2_d, b2_e, b2_v, b2_b, b3_d, b3_e, b3_v, b3_b, b4_d, b4_e, b4_v, b4_b, b5_d, b5_e, b5_v, b5_b, b6_d, b6_e, b6_v, b6_b, b7_d, b7_e, b7_v, b7_b);

  input  clock;
  input  reset;

  input  [15:0] a0_d;
  input  a0_e;
  input  a0_v;
  output a0_b;
  input  [15:0] a1_d;
  input  a1_e;
  input  a1_v;
  output a1_b;
  input  [15:0] a2_d;
  input  a2_e;
  input  a2_v;
  output a2_b;
  input  [15:0] a3_d;
  input  a3_e;
  input  a3_v;
  output a3_b;
  input  [15:0] a4_d;
  input  a4_e;
  input  a4_v;
  output a4_b;
  input  [15:0] a5_d;
  input  a5_e;
  input  a5_v;
  output a5_b;
  input  [15:0] a6_d;
  input  a6_e;
  input  a6_v;
  output a6_b;
  input  [15:0] a7_d;
  input  a7_e;
  input  a7_v;
  output a7_b;
  output [8:0] b0_d;
  output b0_e;
  output b0_v;
  input  b0_b;
  output [8:0] b1_d;
  output b1_e;
  output b1_v;
  input  b1_b;
  output [8:0] b2_d;
  output b2_e;
  output b2_v;
  input  b2_b;
  output [8:0] b3_d;
  output b3_e;
  output b3_v;
  input  b3_b;
  output [8:0] b4_d;
  output b4_e;
  output b4_v;
  input  b4_b;
  output [8:0] b5_d;
  output b5_e;
  output b5_v;
  input  b5_b;
  output [8:0] b6_d;
  output b6_e;
  output b6_v;
  input  b6_b;
  output [8:0] b7_d;
  output b7_e;
  output b7_v;
  input  b7_b;

  wire statecase;

  illm_d1_ScOrEtMp48_fsm fsm (clock, reset, a0_e, a0_v, a0_b, a1_e, a1_v, a1_b, a2_e, a2_v, a2_b, a3_e, a3_v, a3_b, a4_e, a4_v, a4_b, a5_e, a5_v, a5_b, a6_e, a6_v, a6_b, a7_e, a7_v, a7_b, b0_e, b0_v, b0_b, b1_e, b1_v, b1_b, b2_e, b2_v, b2_b, b3_e, b3_v, b3_b, b4_e, b4_v, b4_b, b5_e, b5_v, b5_b, b6_e, b6_v, b6_b, b7_e, b7_v, b7_b, statecase);
  illm_d1_ScOrEtMp48_dp dp (clock, reset, a0_d, a1_d, a2_d, a3_d, a4_d, a5_d, a6_d, a7_d, b0_d, b1_d, b2_d, b3_d, b4_d, b5_d, b6_d, b7_d, statecase);

endmodule  // illm_d1_ScOrEtMp48

module _page_illm_d1_ScOrEtMp48_dpq (clock, reset, a0_d, a0_e, a0_v, a0_b, a1_d, a1_e, a1_v, a1_b, a2_d, a2_e, a2_v, a2_b, a3_d, a3_e, a3_v, a3_b, a4_d, a4_e, a4_v, a4_b, a5_d, a5_e, a5_v, a5_b, a6_d, a6_e, a6_v, a6_b, a7_d, a7_e, a7_v, a7_b, b0_d, b0_e, b0_v, b0_b, b1_d, b1_e, b1_v, b1_b, b2_d, b2_e, b2_v, b2_b, b3_d, b3_e, b3_v, b3_b, b4_d, b4_e, b4_v, b4_b, b5_d, b5_e, b5_v, b5_b, b6_d, b6_e, b6_v, b6_b, b7_d, b7_e, b7_v, b7_b);

  input  clock;
  input  reset;

  input  [15:0] a0_d;
  input  a0_e;
  input  a0_v;
  output a0_b;
  input  [15:0] a1_d;
  input  a1_e;
  input  a1_v;
  output a1_b;
  input  [15:0] a2_d;
  input  a2_e;
  input  a2_v;
  output a2_b;
  input  [15:0] a3_d;
  input  a3_e;
  input  a3_v;
  output a3_b;
  input  [15:0] a4_d;
  input  a4_e;
  input  a4_v;
  output a4_b;
  input  [15:0] a5_d;
  input  a5_e;
  input  a5_v;
  output a5_b;
  input  [15:0] a6_d;
  input  a6_e;
  input  a6_v;
  output a6_b;
  input  [15:0] a7_d;
  input  a7_e;
  input  a7_v;
  output a7_b;
  output [8:0] b0_d;
  output b0_e;
  output b0_v;
  input  b0_b;
  output [8:0] b1_d;
  output b1_e;
  output b1_v;
  input  b1_b;
  output [8:0] b2_d;
  output b2_e;
  output b2_v;
  input  b2_b;
  output [8:0] b3_d;
  output b3_e;
  output b3_v;
  input  b3_b;
  output [8:0] b4_d;
  output b4_e;
  output b4_v;
  input  b4_b;
  output [8:0] b5_d;
  output b5_e;
  output b5_v;
  input  b5_b;
  output [8:0] b6_d;
  output b6_e;
  output b6_v;
  input  b6_b;
  output [8:0] b7_d;
  output b7_e;
  output b7_v;
  input  b7_b;

  wire   [15:0] a0_qin_d, a0_qout_d;
  wire   a0_qin_e, a0_qout_e;
  wire   a0_qin_v, a0_qout_v;
  wire   a0_qin_b, a0_qout_b;
  wire   [15:0] a1_qin_d, a1_qout_d;
  wire   a1_qin_e, a1_qout_e;
  wire   a1_qin_v, a1_qout_v;
  wire   a1_qin_b, a1_qout_b;
  wire   [15:0] a2_qin_d, a2_qout_d;
  wire   a2_qin_e, a2_qout_e;
  wire   a2_qin_v, a2_qout_v;
  wire   a2_qin_b, a2_qout_b;
  wire   [15:0] a3_qin_d, a3_qout_d;
  wire   a3_qin_e, a3_qout_e;
  wire   a3_qin_v, a3_qout_v;
  wire   a3_qin_b, a3_qout_b;
  wire   [15:0] a4_qin_d, a4_qout_d;
  wire   a4_qin_e, a4_qout_e;
  wire   a4_qin_v, a4_qout_v;
  wire   a4_qin_b, a4_qout_b;
  wire   [15:0] a5_qin_d, a5_qout_d;
  wire   a5_qin_e, a5_qout_e;
  wire   a5_qin_v, a5_qout_v;
  wire   a5_qin_b, a5_qout_b;
  wire   [15:0] a6_qin_d, a6_qout_d;
  wire   a6_qin_e, a6_qout_e;
  wire   a6_qin_v, a6_qout_v;
  wire   a6_qin_b, a6_qout_b;
  wire   [15:0] a7_qin_d, a7_qout_d;
  wire   a7_qin_e, a7_qout_e;
  wire   a7_qin_v, a7_qout_v;
  wire   a7_qin_b, a7_qout_b;
  wire   [8:0] b0_qin_d, b0_qout_d;
  wire   b0_qin_e, b0_qout_e;
  wire   b0_qin_v, b0_qout_v;
  wire   b0_qin_b, b0_qout_b;
  wire   [8:0] b1_qin_d, b1_qout_d;
  wire   b1_qin_e, b1_qout_e;
  wire   b1_qin_v, b1_qout_v;
  wire   b1_qin_b, b1_qout_b;
  wire   [8:0] b2_qin_d, b2_qout_d;
  wire   b2_qin_e, b2_qout_e;
  wire   b2_qin_v, b2_qout_v;
  wire   b2_qin_b, b2_qout_b;
  wire   [8:0] b3_qin_d, b3_qout_d;
  wire   b3_qin_e, b3_qout_e;
  wire   b3_qin_v, b3_qout_v;
  wire   b3_qin_b, b3_qout_b;
  wire   [8:0] b4_qin_d, b4_qout_d;
  wire   b4_qin_e, b4_qout_e;
  wire   b4_qin_v, b4_qout_v;
  wire   b4_qin_b, b4_qout_b;
  wire   [8:0] b5_qin_d, b5_qout_d;
  wire   b5_qin_e, b5_qout_e;
  wire   b5_qin_v, b5_qout_v;
  wire   b5_qin_b, b5_qout_b;
  wire   [8:0] b6_qin_d, b6_qout_d;
  wire   b6_qin_e, b6_qout_e;
  wire   b6_qin_v, b6_qout_v;
  wire   b6_qin_b, b6_qout_b;
  wire   [8:0] b7_qin_d, b7_qout_d;
  wire   b7_qin_e, b7_qout_e;
  wire   b7_qin_v, b7_qout_v;
  wire   b7_qin_b, b7_qout_b;

  assign a0_qout_d = a0_d;
  assign a0_qout_e = a0_e;
  assign a0_qout_v = a0_v;
  assign a0_b = a0_qout_b;
  assign a1_qout_d = a1_d;
  assign a1_qout_e = a1_e;
  assign a1_qout_v = a1_v;
  assign a1_b = a1_qout_b;
  assign a2_qout_d = a2_d;
  assign a2_qout_e = a2_e;
  assign a2_qout_v = a2_v;
  assign a2_b = a2_qout_b;
  assign a3_qout_d = a3_d;
  assign a3_qout_e = a3_e;
  assign a3_qout_v = a3_v;
  assign a3_b = a3_qout_b;
  assign a4_qout_d = a4_d;
  assign a4_qout_e = a4_e;
  assign a4_qout_v = a4_v;
  assign a4_b = a4_qout_b;
  assign a5_qout_d = a5_d;
  assign a5_qout_e = a5_e;
  assign a5_qout_v = a5_v;
  assign a5_b = a5_qout_b;
  assign a6_qout_d = a6_d;
  assign a6_qout_e = a6_e;
  assign a6_qout_v = a6_v;
  assign a6_b = a6_qout_b;
  assign a7_qout_d = a7_d;
  assign a7_qout_e = a7_e;
  assign a7_qout_v = a7_v;
  assign a7_b = a7_qout_b;
  assign b0_d = b0_qout_d;
  assign b0_e = b0_qout_e;
  assign b0_v = b0_qout_v;
  assign b0_qout_b = b0_b;
  assign b1_d = b1_qout_d;
  assign b1_e = b1_qout_e;
  assign b1_v = b1_qout_v;
  assign b1_qout_b = b1_b;
  assign b2_d = b2_qout_d;
  assign b2_e = b2_qout_e;
  assign b2_v = b2_qout_v;
  assign b2_qout_b = b2_b;
  assign b3_d = b3_qout_d;
  assign b3_e = b3_qout_e;
  assign b3_v = b3_qout_v;
  assign b3_qout_b = b3_b;
  assign b4_d = b4_qout_d;
  assign b4_e = b4_qout_e;
  assign b4_v = b4_qout_v;
  assign b4_qout_b = b4_b;
  assign b5_d = b5_qout_d;
  assign b5_e = b5_qout_e;
  assign b5_v = b5_qout_v;
  assign b5_qout_b = b5_b;
  assign b6_d = b6_qout_d;
  assign b6_e = b6_qout_e;
  assign b6_v = b6_qout_v;
  assign b6_qout_b = b6_b;
  assign b7_d = b7_qout_d;
  assign b7_e = b7_qout_e;
  assign b7_v = b7_qout_v;
  assign b7_qout_b = b7_b;

  _page_illm_d1_ScOrEtMp48_q _page_illm_d1_ScOrEtMp48_q_ (clock, reset, b0_qin_d, b0_qin_e, b0_qin_v, b0_qin_b, b0_qout_d, b0_qout_e, b0_qout_v, b0_qout_b, b1_qin_d, b1_qin_e, b1_qin_v, b1_qin_b, b1_qout_d, b1_qout_e, b1_qout_v, b1_qout_b, b2_qin_d, b2_qin_e, b2_qin_v, b2_qin_b, b2_qout_d, b2_qout_e, b2_qout_v, b2_qout_b, b3_qin_d, b3_qin_e, b3_qin_v, b3_qin_b, b3_qout_d, b3_qout_e, b3_qout_v, b3_qout_b, b4_qin_d, b4_qin_e, b4_qin_v, b4_qin_b, b4_qout_d, b4_qout_e, b4_qout_v, b4_qout_b, b5_qin_d, b5_qin_e, b5_qin_v, b5_qin_b, b5_qout_d, b5_qout_e, b5_qout_v, b5_qout_b, b6_qin_d, b6_qin_e, b6_qin_v, b6_qin_b, b6_qout_d, b6_qout_e, b6_qout_v, b6_qout_b, b7_qin_d, b7_qin_e, b7_qin_v, b7_qin_b, b7_qout_d, b7_qout_e, b7_qout_v, b7_qout_b);

  illm_d1_ScOrEtMp48 illm_d1_ScOrEtMp48_ (clock, reset, a0_qout_d, a0_qout_e, a0_qout_v, a0_qout_b, a1_qout_d, a1_qout_e, a1_qout_v, a1_qout_b, a2_qout_d, a2_qout_e, a2_qout_v, a2_qout_b, a3_qout_d, a3_qout_e, a3_qout_v, a3_qout_b, a4_qout_d, a4_qout_e, a4_qout_v, a4_qout_b, a5_qout_d, a5_qout_e, a5_qout_v, a5_qout_b, a6_qout_d, a6_qout_e, a6_qout_v, a6_qout_b, a7_qout_d, a7_qout_e, a7_qout_v, a7_qout_b, b0_qin_d, b0_qin_e, b0_qin_v, b0_qin_b, b1_qin_d, b1_qin_e, b1_qin_v, b1_qin_b, b2_qin_d, b2_qin_e, b2_qin_v, b2_qin_b, b3_qin_d, b3_qin_e, b3_qin_v, b3_qin_b, b4_qin_d, b4_qin_e, b4_qin_v, b4_qin_b, b5_qin_d, b5_qin_e, b5_qin_v, b5_qin_b, b6_qin_d, b6_qin_e, b6_qin_v, b6_qin_b, b7_qin_d, b7_qin_e, b7_qin_v, b7_qin_b);

endmodule  // _page_illm_d1_ScOrEtMp48_dpq
