// Verilog inter-page module without input queues for JPEG_dec_d1_ScOrEtMp0
// Emitted by ../../../tdfc version 1.160, Mon Aug 24 17:52:43 2009

`include "JPEG_dec_d1_ScOrEtMp0_q.v"
`include "_page_illm_d1_ScOrEtMp46.v"
`include "_page_tpose_d1_ScOrEtMp47.v"
`include "_page_illm_d1_ScOrEtMp48.v"
`include "_page_bl_d1_ScOrEtMp49.v"
`include "_page_izigzag_d1_ScOrEtMp50.v"
`include "_page_jdquant_d1_ScOrEtMp51.v"
`include "_page_DecHuff_d1_ScOrEtMp52.v"
`include "_page_DecSym_d1_ScOrEtMp53.v"
`include "_page_ftabmod_noinline_d1_ScOrEtMp57.v"
`include "segment_r_0.v"

module JPEG_dec_d1_ScOrEtMp0_noin (clock, reset, outA_d, outA_e, outA_v, outA_b, outB_d, outB_e, outB_v, outB_b, outC_d, outC_e, outC_v, outC_b, outD_d, outD_e, outD_v, outD_b, outE_d, outE_e, outE_v, outE_b, outF_d, outF_e, outF_v, outF_b, outG_d, outG_e, outG_v, outG_b, outH_d, outH_e, outH_v, outH_b, Huffin_d, Huffin_e, Huffin_v, Huffin_b);

  input  clock;
  input  reset;

  output [8:0] outA_d;
  output outA_e;
  output outA_v;
  input  outA_b;
  output [8:0] outB_d;
  output outB_e;
  output outB_v;
  input  outB_b;
  output [8:0] outC_d;
  output outC_e;
  output outC_v;
  input  outC_b;
  output [8:0] outD_d;
  output outD_e;
  output outD_v;
  input  outD_b;
  output [8:0] outE_d;
  output outE_e;
  output outE_v;
  input  outE_b;
  output [8:0] outF_d;
  output outF_e;
  output outF_v;
  input  outF_b;
  output [8:0] outG_d;
  output outG_e;
  output outG_v;
  input  outG_b;
  output [8:0] outH_d;
  output outH_e;
  output outH_v;
  input  outH_b;
  input  [7:0] Huffin_d;
  input  Huffin_e;
  input  Huffin_v;
  output Huffin_b;

  wire   [8:0] outA_qin_d, outA_qout_d;
  wire   outA_qin_e, outA_qout_e;
  wire   outA_qin_v, outA_qout_v;
  wire   outA_qin_b, outA_qout_b;
  wire   [8:0] outB_qin_d, outB_qout_d;
  wire   outB_qin_e, outB_qout_e;
  wire   outB_qin_v, outB_qout_v;
  wire   outB_qin_b, outB_qout_b;
  wire   [8:0] outC_qin_d, outC_qout_d;
  wire   outC_qin_e, outC_qout_e;
  wire   outC_qin_v, outC_qout_v;
  wire   outC_qin_b, outC_qout_b;
  wire   [8:0] outD_qin_d, outD_qout_d;
  wire   outD_qin_e, outD_qout_e;
  wire   outD_qin_v, outD_qout_v;
  wire   outD_qin_b, outD_qout_b;
  wire   [8:0] outE_qin_d, outE_qout_d;
  wire   outE_qin_e, outE_qout_e;
  wire   outE_qin_v, outE_qout_v;
  wire   outE_qin_b, outE_qout_b;
  wire   [8:0] outF_qin_d, outF_qout_d;
  wire   outF_qin_e, outF_qout_e;
  wire   outF_qin_v, outF_qout_v;
  wire   outF_qin_b, outF_qout_b;
  wire   [8:0] outG_qin_d, outG_qout_d;
  wire   outG_qin_e, outG_qout_e;
  wire   outG_qin_v, outG_qout_v;
  wire   outG_qin_b, outG_qout_b;
  wire   [8:0] outH_qin_d, outH_qout_d;
  wire   outH_qin_e, outH_qout_e;
  wire   outH_qin_v, outH_qout_v;
  wire   outH_qin_b, outH_qout_b;
  wire   [7:0] Huffin_qin_d, Huffin_qout_d;
  wire   Huffin_qin_e, Huffin_qout_e;
  wire   Huffin_qin_v, Huffin_qout_v;
  wire   Huffin_qin_b, Huffin_qout_b;
  wire   [15:0] ScOrEtMp1_qin_d, ScOrEtMp1_qout_d;
  wire   ScOrEtMp1_qin_v, ScOrEtMp1_qout_v;
  wire   ScOrEtMp1_qin_e, ScOrEtMp1_qout_e;
  wire   ScOrEtMp1_qin_b, ScOrEtMp1_qout_b;
  wire   [15:0] ScOrEtMp2_qin_d, ScOrEtMp2_qout_d;
  wire   ScOrEtMp2_qin_v, ScOrEtMp2_qout_v;
  wire   ScOrEtMp2_qin_e, ScOrEtMp2_qout_e;
  wire   ScOrEtMp2_qin_b, ScOrEtMp2_qout_b;
  wire   [15:0] ScOrEtMp3_qin_d, ScOrEtMp3_qout_d;
  wire   ScOrEtMp3_qin_v, ScOrEtMp3_qout_v;
  wire   ScOrEtMp3_qin_e, ScOrEtMp3_qout_e;
  wire   ScOrEtMp3_qin_b, ScOrEtMp3_qout_b;
  wire   [15:0] ScOrEtMp4_qin_d, ScOrEtMp4_qout_d;
  wire   ScOrEtMp4_qin_v, ScOrEtMp4_qout_v;
  wire   ScOrEtMp4_qin_e, ScOrEtMp4_qout_e;
  wire   ScOrEtMp4_qin_b, ScOrEtMp4_qout_b;
  wire   [15:0] ScOrEtMp5_qin_d, ScOrEtMp5_qout_d;
  wire   ScOrEtMp5_qin_v, ScOrEtMp5_qout_v;
  wire   ScOrEtMp5_qin_e, ScOrEtMp5_qout_e;
  wire   ScOrEtMp5_qin_b, ScOrEtMp5_qout_b;
  wire   [15:0] ScOrEtMp6_qin_d, ScOrEtMp6_qout_d;
  wire   ScOrEtMp6_qin_v, ScOrEtMp6_qout_v;
  wire   ScOrEtMp6_qin_e, ScOrEtMp6_qout_e;
  wire   ScOrEtMp6_qin_b, ScOrEtMp6_qout_b;
  wire   [15:0] ScOrEtMp7_qin_d, ScOrEtMp7_qout_d;
  wire   ScOrEtMp7_qin_v, ScOrEtMp7_qout_v;
  wire   ScOrEtMp7_qin_e, ScOrEtMp7_qout_e;
  wire   ScOrEtMp7_qin_b, ScOrEtMp7_qout_b;
  wire   [15:0] ScOrEtMp8_qin_d, ScOrEtMp8_qout_d;
  wire   ScOrEtMp8_qin_v, ScOrEtMp8_qout_v;
  wire   ScOrEtMp8_qin_e, ScOrEtMp8_qout_e;
  wire   ScOrEtMp8_qin_b, ScOrEtMp8_qout_b;
  wire   [15:0] ScOrEtMp9_qin_d, ScOrEtMp9_qout_d;
  wire   ScOrEtMp9_qin_v, ScOrEtMp9_qout_v;
  wire   ScOrEtMp9_qin_e, ScOrEtMp9_qout_e;
  wire   ScOrEtMp9_qin_b, ScOrEtMp9_qout_b;
  wire   [15:0] ScOrEtMp10_qin_d, ScOrEtMp10_qout_d;
  wire   ScOrEtMp10_qin_v, ScOrEtMp10_qout_v;
  wire   ScOrEtMp10_qin_e, ScOrEtMp10_qout_e;
  wire   ScOrEtMp10_qin_b, ScOrEtMp10_qout_b;
  wire   [15:0] ScOrEtMp11_qin_d, ScOrEtMp11_qout_d;
  wire   ScOrEtMp11_qin_v, ScOrEtMp11_qout_v;
  wire   ScOrEtMp11_qin_e, ScOrEtMp11_qout_e;
  wire   ScOrEtMp11_qin_b, ScOrEtMp11_qout_b;
  wire   [7:0] ScOrEtMp12_qin_d, ScOrEtMp12_qout_d;
  wire   ScOrEtMp12_qin_v, ScOrEtMp12_qout_v;
  wire   ScOrEtMp12_qin_e, ScOrEtMp12_qout_e;
  wire   ScOrEtMp12_qin_b, ScOrEtMp12_qout_b;
  wire   [7:0] ScOrEtMp13_qin_d, ScOrEtMp13_qout_d;
  wire   ScOrEtMp13_qin_v, ScOrEtMp13_qout_v;
  wire   ScOrEtMp13_qin_e, ScOrEtMp13_qout_e;
  wire   ScOrEtMp13_qin_b, ScOrEtMp13_qout_b;
  wire   [7:0] ScOrEtMp15_qin_d, ScOrEtMp15_qout_d;
  wire   ScOrEtMp15_qin_v, ScOrEtMp15_qout_v;
  wire   ScOrEtMp15_qin_e, ScOrEtMp15_qout_e;
  wire   ScOrEtMp15_qin_b, ScOrEtMp15_qout_b;
  wire   [7:0] ScOrEtMp16_qin_d, ScOrEtMp16_qout_d;
  wire   ScOrEtMp16_qin_v, ScOrEtMp16_qout_v;
  wire   ScOrEtMp16_qin_e, ScOrEtMp16_qout_e;
  wire   ScOrEtMp16_qin_b, ScOrEtMp16_qout_b;
  wire   [15:0] ScOrEtMp21_qin_d, ScOrEtMp21_qout_d;
  wire   ScOrEtMp21_qin_v, ScOrEtMp21_qout_v;
  wire   ScOrEtMp21_qin_e, ScOrEtMp21_qout_e;
  wire   ScOrEtMp21_qin_b, ScOrEtMp21_qout_b;
  wire   [15:0] ScOrEtMp22_qin_d, ScOrEtMp22_qout_d;
  wire   ScOrEtMp22_qin_v, ScOrEtMp22_qout_v;
  wire   ScOrEtMp22_qin_e, ScOrEtMp22_qout_e;
  wire   ScOrEtMp22_qin_b, ScOrEtMp22_qout_b;
  wire   [15:0] ScOrEtMp23_qin_d, ScOrEtMp23_qout_d;
  wire   ScOrEtMp23_qin_v, ScOrEtMp23_qout_v;
  wire   ScOrEtMp23_qin_e, ScOrEtMp23_qout_e;
  wire   ScOrEtMp23_qin_b, ScOrEtMp23_qout_b;
  wire   [15:0] ScOrEtMp24_qin_d, ScOrEtMp24_qout_d;
  wire   ScOrEtMp24_qin_v, ScOrEtMp24_qout_v;
  wire   ScOrEtMp24_qin_e, ScOrEtMp24_qout_e;
  wire   ScOrEtMp24_qin_b, ScOrEtMp24_qout_b;
  wire   [15:0] ScOrEtMp25_qin_d, ScOrEtMp25_qout_d;
  wire   ScOrEtMp25_qin_v, ScOrEtMp25_qout_v;
  wire   ScOrEtMp25_qin_e, ScOrEtMp25_qout_e;
  wire   ScOrEtMp25_qin_b, ScOrEtMp25_qout_b;
  wire   [15:0] ScOrEtMp26_qin_d, ScOrEtMp26_qout_d;
  wire   ScOrEtMp26_qin_v, ScOrEtMp26_qout_v;
  wire   ScOrEtMp26_qin_e, ScOrEtMp26_qout_e;
  wire   ScOrEtMp26_qin_b, ScOrEtMp26_qout_b;
  wire   [15:0] ScOrEtMp27_qin_d, ScOrEtMp27_qout_d;
  wire   ScOrEtMp27_qin_v, ScOrEtMp27_qout_v;
  wire   ScOrEtMp27_qin_e, ScOrEtMp27_qout_e;
  wire   ScOrEtMp27_qin_b, ScOrEtMp27_qout_b;
  wire   [15:0] ScOrEtMp28_qin_d, ScOrEtMp28_qout_d;
  wire   ScOrEtMp28_qin_v, ScOrEtMp28_qout_v;
  wire   ScOrEtMp28_qin_e, ScOrEtMp28_qout_e;
  wire   ScOrEtMp28_qin_b, ScOrEtMp28_qout_b;
  wire   [15:0] ScOrEtMp29_qin_d, ScOrEtMp29_qout_d;
  wire   ScOrEtMp29_qin_v, ScOrEtMp29_qout_v;
  wire   ScOrEtMp29_qin_e, ScOrEtMp29_qout_e;
  wire   ScOrEtMp29_qin_b, ScOrEtMp29_qout_b;
  wire   [15:0] ScOrEtMp30_qin_d, ScOrEtMp30_qout_d;
  wire   ScOrEtMp30_qin_v, ScOrEtMp30_qout_v;
  wire   ScOrEtMp30_qin_e, ScOrEtMp30_qout_e;
  wire   ScOrEtMp30_qin_b, ScOrEtMp30_qout_b;
  wire   [15:0] ScOrEtMp31_qin_d, ScOrEtMp31_qout_d;
  wire   ScOrEtMp31_qin_v, ScOrEtMp31_qout_v;
  wire   ScOrEtMp31_qin_e, ScOrEtMp31_qout_e;
  wire   ScOrEtMp31_qin_b, ScOrEtMp31_qout_b;
  wire   [15:0] ScOrEtMp32_qin_d, ScOrEtMp32_qout_d;
  wire   ScOrEtMp32_qin_v, ScOrEtMp32_qout_v;
  wire   ScOrEtMp32_qin_e, ScOrEtMp32_qout_e;
  wire   ScOrEtMp32_qin_b, ScOrEtMp32_qout_b;
  wire   [15:0] ScOrEtMp33_qin_d, ScOrEtMp33_qout_d;
  wire   ScOrEtMp33_qin_v, ScOrEtMp33_qout_v;
  wire   ScOrEtMp33_qin_e, ScOrEtMp33_qout_e;
  wire   ScOrEtMp33_qin_b, ScOrEtMp33_qout_b;
  wire   [15:0] ScOrEtMp34_qin_d, ScOrEtMp34_qout_d;
  wire   ScOrEtMp34_qin_v, ScOrEtMp34_qout_v;
  wire   ScOrEtMp34_qin_e, ScOrEtMp34_qout_e;
  wire   ScOrEtMp34_qin_b, ScOrEtMp34_qout_b;
  wire   [15:0] ScOrEtMp35_qin_d, ScOrEtMp35_qout_d;
  wire   ScOrEtMp35_qin_v, ScOrEtMp35_qout_v;
  wire   ScOrEtMp35_qin_e, ScOrEtMp35_qout_e;
  wire   ScOrEtMp35_qin_b, ScOrEtMp35_qout_b;
  wire   [15:0] ScOrEtMp36_qin_d, ScOrEtMp36_qout_d;
  wire   ScOrEtMp36_qin_v, ScOrEtMp36_qout_v;
  wire   ScOrEtMp36_qin_e, ScOrEtMp36_qout_e;
  wire   ScOrEtMp36_qin_b, ScOrEtMp36_qout_b;
  wire   [8:0] ScOrEtMp37_qin_d, ScOrEtMp37_qout_d;
  wire   ScOrEtMp37_qin_v, ScOrEtMp37_qout_v;
  wire   ScOrEtMp37_qin_e, ScOrEtMp37_qout_e;
  wire   ScOrEtMp37_qin_b, ScOrEtMp37_qout_b;
  wire   [8:0] ScOrEtMp38_qin_d, ScOrEtMp38_qout_d;
  wire   ScOrEtMp38_qin_v, ScOrEtMp38_qout_v;
  wire   ScOrEtMp38_qin_e, ScOrEtMp38_qout_e;
  wire   ScOrEtMp38_qin_b, ScOrEtMp38_qout_b;
  wire   [8:0] ScOrEtMp39_qin_d, ScOrEtMp39_qout_d;
  wire   ScOrEtMp39_qin_v, ScOrEtMp39_qout_v;
  wire   ScOrEtMp39_qin_e, ScOrEtMp39_qout_e;
  wire   ScOrEtMp39_qin_b, ScOrEtMp39_qout_b;
  wire   [8:0] ScOrEtMp40_qin_d, ScOrEtMp40_qout_d;
  wire   ScOrEtMp40_qin_v, ScOrEtMp40_qout_v;
  wire   ScOrEtMp40_qin_e, ScOrEtMp40_qout_e;
  wire   ScOrEtMp40_qin_b, ScOrEtMp40_qout_b;
  wire   [8:0] ScOrEtMp41_qin_d, ScOrEtMp41_qout_d;
  wire   ScOrEtMp41_qin_v, ScOrEtMp41_qout_v;
  wire   ScOrEtMp41_qin_e, ScOrEtMp41_qout_e;
  wire   ScOrEtMp41_qin_b, ScOrEtMp41_qout_b;
  wire   [8:0] ScOrEtMp42_qin_d, ScOrEtMp42_qout_d;
  wire   ScOrEtMp42_qin_v, ScOrEtMp42_qout_v;
  wire   ScOrEtMp42_qin_e, ScOrEtMp42_qout_e;
  wire   ScOrEtMp42_qin_b, ScOrEtMp42_qout_b;
  wire   [8:0] ScOrEtMp43_qin_d, ScOrEtMp43_qout_d;
  wire   ScOrEtMp43_qin_v, ScOrEtMp43_qout_v;
  wire   ScOrEtMp43_qin_e, ScOrEtMp43_qout_e;
  wire   ScOrEtMp43_qin_b, ScOrEtMp43_qout_b;
  wire   [8:0] ScOrEtMp44_qin_d, ScOrEtMp44_qout_d;
  wire   ScOrEtMp44_qin_v, ScOrEtMp44_qout_v;
  wire   ScOrEtMp44_qin_e, ScOrEtMp44_qout_e;
  wire   ScOrEtMp44_qin_b, ScOrEtMp44_qout_b;
  wire   [31:0] ScOrEtMp55_qin_d, ScOrEtMp55_qout_d;
  wire   ScOrEtMp55_qin_v, ScOrEtMp55_qout_v;
  wire   ScOrEtMp55_qin_e, ScOrEtMp55_qout_e;
  wire   ScOrEtMp55_qin_b, ScOrEtMp55_qout_b;
  wire   [63:0] ScOrEtMp56_qin_d, ScOrEtMp56_qout_d;
  wire   ScOrEtMp56_qin_v, ScOrEtMp56_qout_v;
  wire   ScOrEtMp56_qin_e, ScOrEtMp56_qout_e;
  wire   ScOrEtMp56_qin_b, ScOrEtMp56_qout_b;

  assign outA_d = outA_qout_d;
  assign outA_e = outA_qout_e;
  assign outA_v = outA_qout_v;
  assign outA_qout_b = outA_b;
  assign outB_d = outB_qout_d;
  assign outB_e = outB_qout_e;
  assign outB_v = outB_qout_v;
  assign outB_qout_b = outB_b;
  assign outC_d = outC_qout_d;
  assign outC_e = outC_qout_e;
  assign outC_v = outC_qout_v;
  assign outC_qout_b = outC_b;
  assign outD_d = outD_qout_d;
  assign outD_e = outD_qout_e;
  assign outD_v = outD_qout_v;
  assign outD_qout_b = outD_b;
  assign outE_d = outE_qout_d;
  assign outE_e = outE_qout_e;
  assign outE_v = outE_qout_v;
  assign outE_qout_b = outE_b;
  assign outF_d = outF_qout_d;
  assign outF_e = outF_qout_e;
  assign outF_v = outF_qout_v;
  assign outF_qout_b = outF_b;
  assign outG_d = outG_qout_d;
  assign outG_e = outG_qout_e;
  assign outG_v = outG_qout_v;
  assign outG_qout_b = outG_b;
  assign outH_d = outH_qout_d;
  assign outH_e = outH_qout_e;
  assign outH_v = outH_qout_v;
  assign outH_qout_b = outH_b;
  assign Huffin_qout_d = Huffin_d;
  assign Huffin_qout_e = Huffin_e;
  assign Huffin_qout_v = Huffin_v;
  assign Huffin_b = Huffin_qout_b;

  JPEG_dec_d1_ScOrEtMp0_q JPEG_dec_d1_ScOrEtMp0_q_ (clock, reset, outA_qin_d, outA_qin_e, outA_qin_v, outA_qin_b, outA_qout_d, outA_qout_e, outA_qout_v, outA_qout_b, outB_qin_d, outB_qin_e, outB_qin_v, outB_qin_b, outB_qout_d, outB_qout_e, outB_qout_v, outB_qout_b, outC_qin_d, outC_qin_e, outC_qin_v, outC_qin_b, outC_qout_d, outC_qout_e, outC_qout_v, outC_qout_b, outD_qin_d, outD_qin_e, outD_qin_v, outD_qin_b, outD_qout_d, outD_qout_e, outD_qout_v, outD_qout_b, outE_qin_d, outE_qin_e, outE_qin_v, outE_qin_b, outE_qout_d, outE_qout_e, outE_qout_v, outE_qout_b, outF_qin_d, outF_qin_e, outF_qin_v, outF_qin_b, outF_qout_d, outF_qout_e, outF_qout_v, outF_qout_b, outG_qin_d, outG_qin_e, outG_qin_v, outG_qin_b, outG_qout_d, outG_qout_e, outG_qout_v, outG_qout_b, outH_qin_d, outH_qin_e, outH_qin_v, outH_qin_b, outH_qout_d, outH_qout_e, outH_qout_v, outH_qout_b, ScOrEtMp1_qin_d, ScOrEtMp1_qin_e, ScOrEtMp1_qin_v, ScOrEtMp1_qin_b, ScOrEtMp1_qout_d, ScOrEtMp1_qout_e, ScOrEtMp1_qout_v, ScOrEtMp1_qout_b, ScOrEtMp2_qin_d, ScOrEtMp2_qin_e, ScOrEtMp2_qin_v, ScOrEtMp2_qin_b, ScOrEtMp2_qout_d, ScOrEtMp2_qout_e, ScOrEtMp2_qout_v, ScOrEtMp2_qout_b, ScOrEtMp3_qin_d, ScOrEtMp3_qin_e, ScOrEtMp3_qin_v, ScOrEtMp3_qin_b, ScOrEtMp3_qout_d, ScOrEtMp3_qout_e, ScOrEtMp3_qout_v, ScOrEtMp3_qout_b, ScOrEtMp4_qin_d, ScOrEtMp4_qin_e, ScOrEtMp4_qin_v, ScOrEtMp4_qin_b, ScOrEtMp4_qout_d, ScOrEtMp4_qout_e, ScOrEtMp4_qout_v, ScOrEtMp4_qout_b, ScOrEtMp5_qin_d, ScOrEtMp5_qin_e, ScOrEtMp5_qin_v, ScOrEtMp5_qin_b, ScOrEtMp5_qout_d, ScOrEtMp5_qout_e, ScOrEtMp5_qout_v, ScOrEtMp5_qout_b, ScOrEtMp6_qin_d, ScOrEtMp6_qin_e, ScOrEtMp6_qin_v, ScOrEtMp6_qin_b, ScOrEtMp6_qout_d, ScOrEtMp6_qout_e, ScOrEtMp6_qout_v, ScOrEtMp6_qout_b, ScOrEtMp7_qin_d, ScOrEtMp7_qin_e, ScOrEtMp7_qin_v, ScOrEtMp7_qin_b, ScOrEtMp7_qout_d, ScOrEtMp7_qout_e, ScOrEtMp7_qout_v, ScOrEtMp7_qout_b, ScOrEtMp8_qin_d, ScOrEtMp8_qin_e, ScOrEtMp8_qin_v, ScOrEtMp8_qin_b, ScOrEtMp8_qout_d, ScOrEtMp8_qout_e, ScOrEtMp8_qout_v, ScOrEtMp8_qout_b, ScOrEtMp9_qin_d, ScOrEtMp9_qin_e, ScOrEtMp9_qin_v, ScOrEtMp9_qin_b, ScOrEtMp9_qout_d, ScOrEtMp9_qout_e, ScOrEtMp9_qout_v, ScOrEtMp9_qout_b, ScOrEtMp10_qin_d, ScOrEtMp10_qin_e, ScOrEtMp10_qin_v, ScOrEtMp10_qin_b, ScOrEtMp10_qout_d, ScOrEtMp10_qout_e, ScOrEtMp10_qout_v, ScOrEtMp10_qout_b, ScOrEtMp11_qin_d, ScOrEtMp11_qin_e, ScOrEtMp11_qin_v, ScOrEtMp11_qin_b, ScOrEtMp11_qout_d, ScOrEtMp11_qout_e, ScOrEtMp11_qout_v, ScOrEtMp11_qout_b, ScOrEtMp12_qin_d, ScOrEtMp12_qin_e, ScOrEtMp12_qin_v, ScOrEtMp12_qin_b, ScOrEtMp12_qout_d, ScOrEtMp12_qout_e, ScOrEtMp12_qout_v, ScOrEtMp12_qout_b, ScOrEtMp13_qin_d, ScOrEtMp13_qin_e, ScOrEtMp13_qin_v, ScOrEtMp13_qin_b, ScOrEtMp13_qout_d, ScOrEtMp13_qout_e, ScOrEtMp13_qout_v, ScOrEtMp13_qout_b, ScOrEtMp15_qin_d, ScOrEtMp15_qin_e, ScOrEtMp15_qin_v, ScOrEtMp15_qin_b, ScOrEtMp15_qout_d, ScOrEtMp15_qout_e, ScOrEtMp15_qout_v, ScOrEtMp15_qout_b, ScOrEtMp16_qin_d, ScOrEtMp16_qin_e, ScOrEtMp16_qin_v, ScOrEtMp16_qin_b, ScOrEtMp16_qout_d, ScOrEtMp16_qout_e, ScOrEtMp16_qout_v, ScOrEtMp16_qout_b, ScOrEtMp21_qin_d, ScOrEtMp21_qin_e, ScOrEtMp21_qin_v, ScOrEtMp21_qin_b, ScOrEtMp21_qout_d, ScOrEtMp21_qout_e, ScOrEtMp21_qout_v, ScOrEtMp21_qout_b, ScOrEtMp22_qin_d, ScOrEtMp22_qin_e, ScOrEtMp22_qin_v, ScOrEtMp22_qin_b, ScOrEtMp22_qout_d, ScOrEtMp22_qout_e, ScOrEtMp22_qout_v, ScOrEtMp22_qout_b, ScOrEtMp23_qin_d, ScOrEtMp23_qin_e, ScOrEtMp23_qin_v, ScOrEtMp23_qin_b, ScOrEtMp23_qout_d, ScOrEtMp23_qout_e, ScOrEtMp23_qout_v, ScOrEtMp23_qout_b, ScOrEtMp24_qin_d, ScOrEtMp24_qin_e, ScOrEtMp24_qin_v, ScOrEtMp24_qin_b, ScOrEtMp24_qout_d, ScOrEtMp24_qout_e, ScOrEtMp24_qout_v, ScOrEtMp24_qout_b, ScOrEtMp25_qin_d, ScOrEtMp25_qin_e, ScOrEtMp25_qin_v, ScOrEtMp25_qin_b, ScOrEtMp25_qout_d, ScOrEtMp25_qout_e, ScOrEtMp25_qout_v, ScOrEtMp25_qout_b, ScOrEtMp26_qin_d, ScOrEtMp26_qin_e, ScOrEtMp26_qin_v, ScOrEtMp26_qin_b, ScOrEtMp26_qout_d, ScOrEtMp26_qout_e, ScOrEtMp26_qout_v, ScOrEtMp26_qout_b, ScOrEtMp27_qin_d, ScOrEtMp27_qin_e, ScOrEtMp27_qin_v, ScOrEtMp27_qin_b, ScOrEtMp27_qout_d, ScOrEtMp27_qout_e, ScOrEtMp27_qout_v, ScOrEtMp27_qout_b, ScOrEtMp28_qin_d, ScOrEtMp28_qin_e, ScOrEtMp28_qin_v, ScOrEtMp28_qin_b, ScOrEtMp28_qout_d, ScOrEtMp28_qout_e, ScOrEtMp28_qout_v, ScOrEtMp28_qout_b, ScOrEtMp29_qin_d, ScOrEtMp29_qin_e, ScOrEtMp29_qin_v, ScOrEtMp29_qin_b, ScOrEtMp29_qout_d, ScOrEtMp29_qout_e, ScOrEtMp29_qout_v, ScOrEtMp29_qout_b, ScOrEtMp30_qin_d, ScOrEtMp30_qin_e, ScOrEtMp30_qin_v, ScOrEtMp30_qin_b, ScOrEtMp30_qout_d, ScOrEtMp30_qout_e, ScOrEtMp30_qout_v, ScOrEtMp30_qout_b, ScOrEtMp31_qin_d, ScOrEtMp31_qin_e, ScOrEtMp31_qin_v, ScOrEtMp31_qin_b, ScOrEtMp31_qout_d, ScOrEtMp31_qout_e, ScOrEtMp31_qout_v, ScOrEtMp31_qout_b, ScOrEtMp32_qin_d, ScOrEtMp32_qin_e, ScOrEtMp32_qin_v, ScOrEtMp32_qin_b, ScOrEtMp32_qout_d, ScOrEtMp32_qout_e, ScOrEtMp32_qout_v, ScOrEtMp32_qout_b, ScOrEtMp33_qin_d, ScOrEtMp33_qin_e, ScOrEtMp33_qin_v, ScOrEtMp33_qin_b, ScOrEtMp33_qout_d, ScOrEtMp33_qout_e, ScOrEtMp33_qout_v, ScOrEtMp33_qout_b, ScOrEtMp34_qin_d, ScOrEtMp34_qin_e, ScOrEtMp34_qin_v, ScOrEtMp34_qin_b, ScOrEtMp34_qout_d, ScOrEtMp34_qout_e, ScOrEtMp34_qout_v, ScOrEtMp34_qout_b, ScOrEtMp35_qin_d, ScOrEtMp35_qin_e, ScOrEtMp35_qin_v, ScOrEtMp35_qin_b, ScOrEtMp35_qout_d, ScOrEtMp35_qout_e, ScOrEtMp35_qout_v, ScOrEtMp35_qout_b, ScOrEtMp36_qin_d, ScOrEtMp36_qin_e, ScOrEtMp36_qin_v, ScOrEtMp36_qin_b, ScOrEtMp36_qout_d, ScOrEtMp36_qout_e, ScOrEtMp36_qout_v, ScOrEtMp36_qout_b, ScOrEtMp37_qin_d, ScOrEtMp37_qin_e, ScOrEtMp37_qin_v, ScOrEtMp37_qin_b, ScOrEtMp37_qout_d, ScOrEtMp37_qout_e, ScOrEtMp37_qout_v, ScOrEtMp37_qout_b, ScOrEtMp38_qin_d, ScOrEtMp38_qin_e, ScOrEtMp38_qin_v, ScOrEtMp38_qin_b, ScOrEtMp38_qout_d, ScOrEtMp38_qout_e, ScOrEtMp38_qout_v, ScOrEtMp38_qout_b, ScOrEtMp39_qin_d, ScOrEtMp39_qin_e, ScOrEtMp39_qin_v, ScOrEtMp39_qin_b, ScOrEtMp39_qout_d, ScOrEtMp39_qout_e, ScOrEtMp39_qout_v, ScOrEtMp39_qout_b, ScOrEtMp40_qin_d, ScOrEtMp40_qin_e, ScOrEtMp40_qin_v, ScOrEtMp40_qin_b, ScOrEtMp40_qout_d, ScOrEtMp40_qout_e, ScOrEtMp40_qout_v, ScOrEtMp40_qout_b, ScOrEtMp41_qin_d, ScOrEtMp41_qin_e, ScOrEtMp41_qin_v, ScOrEtMp41_qin_b, ScOrEtMp41_qout_d, ScOrEtMp41_qout_e, ScOrEtMp41_qout_v, ScOrEtMp41_qout_b, ScOrEtMp42_qin_d, ScOrEtMp42_qin_e, ScOrEtMp42_qin_v, ScOrEtMp42_qin_b, ScOrEtMp42_qout_d, ScOrEtMp42_qout_e, ScOrEtMp42_qout_v, ScOrEtMp42_qout_b, ScOrEtMp43_qin_d, ScOrEtMp43_qin_e, ScOrEtMp43_qin_v, ScOrEtMp43_qin_b, ScOrEtMp43_qout_d, ScOrEtMp43_qout_e, ScOrEtMp43_qout_v, ScOrEtMp43_qout_b, ScOrEtMp44_qin_d, ScOrEtMp44_qin_e, ScOrEtMp44_qin_v, ScOrEtMp44_qin_b, ScOrEtMp44_qout_d, ScOrEtMp44_qout_e, ScOrEtMp44_qout_v, ScOrEtMp44_qout_b, ScOrEtMp55_qin_d, ScOrEtMp55_qin_e, ScOrEtMp55_qin_v, ScOrEtMp55_qin_b, ScOrEtMp55_qout_d, ScOrEtMp55_qout_e, ScOrEtMp55_qout_v, ScOrEtMp55_qout_b, ScOrEtMp56_qin_d, ScOrEtMp56_qin_e, ScOrEtMp56_qin_v, ScOrEtMp56_qin_b, ScOrEtMp56_qout_d, ScOrEtMp56_qout_e, ScOrEtMp56_qout_v, ScOrEtMp56_qout_b);

  _page_illm_d1_ScOrEtMp46 _page_illm_d1_ScOrEtMp46_ (clock, reset, ScOrEtMp1_qout_d, ScOrEtMp1_qout_e, ScOrEtMp1_qout_v, ScOrEtMp1_qout_b, ScOrEtMp2_qout_d, ScOrEtMp2_qout_e, ScOrEtMp2_qout_v, ScOrEtMp2_qout_b, ScOrEtMp3_qout_d, ScOrEtMp3_qout_e, ScOrEtMp3_qout_v, ScOrEtMp3_qout_b, ScOrEtMp4_qout_d, ScOrEtMp4_qout_e, ScOrEtMp4_qout_v, ScOrEtMp4_qout_b, ScOrEtMp5_qout_d, ScOrEtMp5_qout_e, ScOrEtMp5_qout_v, ScOrEtMp5_qout_b, ScOrEtMp6_qout_d, ScOrEtMp6_qout_e, ScOrEtMp6_qout_v, ScOrEtMp6_qout_b, ScOrEtMp7_qout_d, ScOrEtMp7_qout_e, ScOrEtMp7_qout_v, ScOrEtMp7_qout_b, ScOrEtMp8_qout_d, ScOrEtMp8_qout_e, ScOrEtMp8_qout_v, ScOrEtMp8_qout_b, ScOrEtMp21_qin_d, ScOrEtMp21_qin_e, ScOrEtMp21_qin_v, ScOrEtMp21_qin_b, ScOrEtMp22_qin_d, ScOrEtMp22_qin_e, ScOrEtMp22_qin_v, ScOrEtMp22_qin_b, ScOrEtMp23_qin_d, ScOrEtMp23_qin_e, ScOrEtMp23_qin_v, ScOrEtMp23_qin_b, ScOrEtMp24_qin_d, ScOrEtMp24_qin_e, ScOrEtMp24_qin_v, ScOrEtMp24_qin_b, ScOrEtMp25_qin_d, ScOrEtMp25_qin_e, ScOrEtMp25_qin_v, ScOrEtMp25_qin_b, ScOrEtMp26_qin_d, ScOrEtMp26_qin_e, ScOrEtMp26_qin_v, ScOrEtMp26_qin_b, ScOrEtMp27_qin_d, ScOrEtMp27_qin_e, ScOrEtMp27_qin_v, ScOrEtMp27_qin_b, ScOrEtMp28_qin_d, ScOrEtMp28_qin_e, ScOrEtMp28_qin_v, ScOrEtMp28_qin_b);
  _page_tpose_d1_ScOrEtMp47 _page_tpose_d1_ScOrEtMp47_ (clock, reset, ScOrEtMp21_qout_d, ScOrEtMp21_qout_e, ScOrEtMp21_qout_v, ScOrEtMp21_qout_b, ScOrEtMp22_qout_d, ScOrEtMp22_qout_e, ScOrEtMp22_qout_v, ScOrEtMp22_qout_b, ScOrEtMp23_qout_d, ScOrEtMp23_qout_e, ScOrEtMp23_qout_v, ScOrEtMp23_qout_b, ScOrEtMp24_qout_d, ScOrEtMp24_qout_e, ScOrEtMp24_qout_v, ScOrEtMp24_qout_b, ScOrEtMp25_qout_d, ScOrEtMp25_qout_e, ScOrEtMp25_qout_v, ScOrEtMp25_qout_b, ScOrEtMp26_qout_d, ScOrEtMp26_qout_e, ScOrEtMp26_qout_v, ScOrEtMp26_qout_b, ScOrEtMp27_qout_d, ScOrEtMp27_qout_e, ScOrEtMp27_qout_v, ScOrEtMp27_qout_b, ScOrEtMp28_qout_d, ScOrEtMp28_qout_e, ScOrEtMp28_qout_v, ScOrEtMp28_qout_b, ScOrEtMp29_qin_d, ScOrEtMp29_qin_e, ScOrEtMp29_qin_v, ScOrEtMp29_qin_b, ScOrEtMp30_qin_d, ScOrEtMp30_qin_e, ScOrEtMp30_qin_v, ScOrEtMp30_qin_b, ScOrEtMp31_qin_d, ScOrEtMp31_qin_e, ScOrEtMp31_qin_v, ScOrEtMp31_qin_b, ScOrEtMp32_qin_d, ScOrEtMp32_qin_e, ScOrEtMp32_qin_v, ScOrEtMp32_qin_b, ScOrEtMp33_qin_d, ScOrEtMp33_qin_e, ScOrEtMp33_qin_v, ScOrEtMp33_qin_b, ScOrEtMp34_qin_d, ScOrEtMp34_qin_e, ScOrEtMp34_qin_v, ScOrEtMp34_qin_b, ScOrEtMp35_qin_d, ScOrEtMp35_qin_e, ScOrEtMp35_qin_v, ScOrEtMp35_qin_b, ScOrEtMp36_qin_d, ScOrEtMp36_qin_e, ScOrEtMp36_qin_v, ScOrEtMp36_qin_b);
  _page_illm_d1_ScOrEtMp48 _page_illm_d1_ScOrEtMp48_ (clock, reset, ScOrEtMp29_qout_d, ScOrEtMp29_qout_e, ScOrEtMp29_qout_v, ScOrEtMp29_qout_b, ScOrEtMp30_qout_d, ScOrEtMp30_qout_e, ScOrEtMp30_qout_v, ScOrEtMp30_qout_b, ScOrEtMp31_qout_d, ScOrEtMp31_qout_e, ScOrEtMp31_qout_v, ScOrEtMp31_qout_b, ScOrEtMp32_qout_d, ScOrEtMp32_qout_e, ScOrEtMp32_qout_v, ScOrEtMp32_qout_b, ScOrEtMp33_qout_d, ScOrEtMp33_qout_e, ScOrEtMp33_qout_v, ScOrEtMp33_qout_b, ScOrEtMp34_qout_d, ScOrEtMp34_qout_e, ScOrEtMp34_qout_v, ScOrEtMp34_qout_b, ScOrEtMp35_qout_d, ScOrEtMp35_qout_e, ScOrEtMp35_qout_v, ScOrEtMp35_qout_b, ScOrEtMp36_qout_d, ScOrEtMp36_qout_e, ScOrEtMp36_qout_v, ScOrEtMp36_qout_b, ScOrEtMp37_qin_d, ScOrEtMp37_qin_e, ScOrEtMp37_qin_v, ScOrEtMp37_qin_b, ScOrEtMp38_qin_d, ScOrEtMp38_qin_e, ScOrEtMp38_qin_v, ScOrEtMp38_qin_b, ScOrEtMp39_qin_d, ScOrEtMp39_qin_e, ScOrEtMp39_qin_v, ScOrEtMp39_qin_b, ScOrEtMp40_qin_d, ScOrEtMp40_qin_e, ScOrEtMp40_qin_v, ScOrEtMp40_qin_b, ScOrEtMp41_qin_d, ScOrEtMp41_qin_e, ScOrEtMp41_qin_v, ScOrEtMp41_qin_b, ScOrEtMp42_qin_d, ScOrEtMp42_qin_e, ScOrEtMp42_qin_v, ScOrEtMp42_qin_b, ScOrEtMp43_qin_d, ScOrEtMp43_qin_e, ScOrEtMp43_qin_v, ScOrEtMp43_qin_b, ScOrEtMp44_qin_d, ScOrEtMp44_qin_e, ScOrEtMp44_qin_v, ScOrEtMp44_qin_b);
  _page_bl_d1_ScOrEtMp49 _page_bl_d1_ScOrEtMp49_ (clock, reset, ScOrEtMp37_qout_d, ScOrEtMp37_qout_e, ScOrEtMp37_qout_v, ScOrEtMp37_qout_b, ScOrEtMp38_qout_d, ScOrEtMp38_qout_e, ScOrEtMp38_qout_v, ScOrEtMp38_qout_b, ScOrEtMp39_qout_d, ScOrEtMp39_qout_e, ScOrEtMp39_qout_v, ScOrEtMp39_qout_b, ScOrEtMp40_qout_d, ScOrEtMp40_qout_e, ScOrEtMp40_qout_v, ScOrEtMp40_qout_b, ScOrEtMp41_qout_d, ScOrEtMp41_qout_e, ScOrEtMp41_qout_v, ScOrEtMp41_qout_b, ScOrEtMp42_qout_d, ScOrEtMp42_qout_e, ScOrEtMp42_qout_v, ScOrEtMp42_qout_b, ScOrEtMp43_qout_d, ScOrEtMp43_qout_e, ScOrEtMp43_qout_v, ScOrEtMp43_qout_b, ScOrEtMp44_qout_d, ScOrEtMp44_qout_e, ScOrEtMp44_qout_v, ScOrEtMp44_qout_b, outA_qin_d, outA_qin_e, outA_qin_v, outA_qin_b, outB_qin_d, outB_qin_e, outB_qin_v, outB_qin_b, outC_qin_d, outC_qin_e, outC_qin_v, outC_qin_b, outD_qin_d, outD_qin_e, outD_qin_v, outD_qin_b, outE_qin_d, outE_qin_e, outE_qin_v, outE_qin_b, outF_qin_d, outF_qin_e, outF_qin_v, outF_qin_b, outG_qin_d, outG_qin_e, outG_qin_v, outG_qin_b, outH_qin_d, outH_qin_e, outH_qin_v, outH_qin_b);
  _page_izigzag_d1_ScOrEtMp50 _page_izigzag_d1_ScOrEtMp50_ (clock, reset, ScOrEtMp1_qin_d, ScOrEtMp1_qin_e, ScOrEtMp1_qin_v, ScOrEtMp1_qin_b, ScOrEtMp2_qin_d, ScOrEtMp2_qin_e, ScOrEtMp2_qin_v, ScOrEtMp2_qin_b, ScOrEtMp3_qin_d, ScOrEtMp3_qin_e, ScOrEtMp3_qin_v, ScOrEtMp3_qin_b, ScOrEtMp4_qin_d, ScOrEtMp4_qin_e, ScOrEtMp4_qin_v, ScOrEtMp4_qin_b, ScOrEtMp5_qin_d, ScOrEtMp5_qin_e, ScOrEtMp5_qin_v, ScOrEtMp5_qin_b, ScOrEtMp6_qin_d, ScOrEtMp6_qin_e, ScOrEtMp6_qin_v, ScOrEtMp6_qin_b, ScOrEtMp7_qin_d, ScOrEtMp7_qin_e, ScOrEtMp7_qin_v, ScOrEtMp7_qin_b, ScOrEtMp8_qin_d, ScOrEtMp8_qin_e, ScOrEtMp8_qin_v, ScOrEtMp8_qin_b, ScOrEtMp9_qout_d, ScOrEtMp9_qout_e, ScOrEtMp9_qout_v, ScOrEtMp9_qout_b);
  _page_jdquant_d1_ScOrEtMp51 _page_jdquant_d1_ScOrEtMp51_ (clock, reset, ScOrEtMp10_qout_d, ScOrEtMp10_qout_e, ScOrEtMp10_qout_v, ScOrEtMp10_qout_b, ScOrEtMp9_qin_d, ScOrEtMp9_qin_e, ScOrEtMp9_qin_v, ScOrEtMp9_qin_b);
  _page_DecHuff_d1_ScOrEtMp52 _page_DecHuff_d1_ScOrEtMp52_ (clock, reset, Huffin_qout_d, Huffin_qout_e, Huffin_qout_v, Huffin_qout_b, ScOrEtMp12_qout_d, ScOrEtMp12_qout_e, ScOrEtMp12_qout_v, ScOrEtMp12_qout_b, ScOrEtMp13_qout_d, ScOrEtMp13_qout_e, ScOrEtMp13_qout_v, ScOrEtMp13_qout_b, ScOrEtMp11_qin_d, ScOrEtMp11_qin_e, ScOrEtMp11_qin_v, ScOrEtMp11_qin_b);
  _page_DecSym_d1_ScOrEtMp53 _page_DecSym_d1_ScOrEtMp53_ (clock, reset, ScOrEtMp11_qout_d, ScOrEtMp11_qout_e, ScOrEtMp11_qout_v, ScOrEtMp11_qout_b, ScOrEtMp13_qin_d, ScOrEtMp13_qin_e, ScOrEtMp13_qin_v, ScOrEtMp13_qin_b, ScOrEtMp12_qin_d, ScOrEtMp12_qin_e, ScOrEtMp12_qin_v, ScOrEtMp12_qin_b, ScOrEtMp10_qin_d, ScOrEtMp10_qin_e, ScOrEtMp10_qin_v, ScOrEtMp10_qin_b, ScOrEtMp15_qin_d, ScOrEtMp15_qin_e, ScOrEtMp15_qin_v, ScOrEtMp15_qin_b, ScOrEtMp16_qout_d, ScOrEtMp16_qout_e, ScOrEtMp16_qout_v, ScOrEtMp16_qout_b);
  _page_ftabmod_noinline_d1_ScOrEtMp57 _page_ftabmod_noinline_d1_ScOrEtMp57_ (clock, reset, ScOrEtMp15_qout_d, ScOrEtMp15_qout_e, ScOrEtMp15_qout_v, ScOrEtMp15_qout_b, ScOrEtMp16_qin_d, ScOrEtMp16_qin_e, ScOrEtMp16_qin_v, ScOrEtMp16_qin_b, ScOrEtMp55_qin_d, ScOrEtMp55_qin_e, ScOrEtMp55_qin_v, ScOrEtMp55_qin_b, ScOrEtMp56_qout_d, ScOrEtMp56_qout_e, ScOrEtMp56_qout_v, ScOrEtMp56_qout_b);
  segment_r_0 segment_r_0_ (clock, reset, ScOrEtMp55_qout_d, ScOrEtMp55_qout_e, ScOrEtMp55_qout_v, ScOrEtMp55_qout_b, ScOrEtMp56_qin_d, ScOrEtMp56_qin_e, ScOrEtMp56_qin_v, ScOrEtMp56_qin_b);

endmodule  // JPEG_dec_d1_ScOrEtMp0_noin
